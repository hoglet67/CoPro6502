library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tuberom_68000 is
    port (
        CLK  : in  std_logic;
        ADDR : in  std_logic_vector(13 downto 0);
        DATA : out std_logic_vector(15 downto 0)
        );
end;

architecture RTL of tuberom_68000 is

    signal rom_addr : std_logic_vector(13 downto 0);

begin

    p_addr : process(ADDR)
    begin
        rom_addr              <= (others => '0');
        rom_addr(13 downto 0) <= ADDR;
    end process;

    p_rom : process
    begin
        wait until rising_edge(CLK);
        DATA <= (others => '0');
        case rom_addr is
            when "00" & x"000" => DATA <= x"0000";
            when "00" & x"001" => DATA <= x"0620";
            when "00" & x"002" => DATA <= x"003f";
            when "00" & x"003" => DATA <= x"0200";
            when "00" & x"004" => DATA <= x"003f";
            when "00" & x"005" => DATA <= x"0626";
            when "00" & x"006" => DATA <= x"003f";
            when "00" & x"007" => DATA <= x"072e";
            when "00" & x"008" => DATA <= x"003f";
            when "00" & x"009" => DATA <= x"073c";
            when "00" & x"00a" => DATA <= x"003f";
            when "00" & x"00b" => DATA <= x"0748";
            when "00" & x"00c" => DATA <= x"003f";
            when "00" & x"00d" => DATA <= x"0760";
            when "00" & x"00e" => DATA <= x"003f";
            when "00" & x"00f" => DATA <= x"0760";
            when "00" & x"010" => DATA <= x"003f";
            when "00" & x"011" => DATA <= x"0754";
            when "00" & x"012" => DATA <= x"003f";
            when "00" & x"013" => DATA <= x"0760";
            when "00" & x"014" => DATA <= x"003f";
            when "00" & x"015" => DATA <= x"0760";
            when "00" & x"016" => DATA <= x"003f";
            when "00" & x"017" => DATA <= x"0760";
            when "00" & x"018" => DATA <= x"003f";
            when "00" & x"019" => DATA <= x"0760";
            when "00" & x"01a" => DATA <= x"003f";
            when "00" & x"01b" => DATA <= x"0760";
            when "00" & x"01c" => DATA <= x"003f";
            when "00" & x"01d" => DATA <= x"0760";
            when "00" & x"01e" => DATA <= x"003f";
            when "00" & x"01f" => DATA <= x"0760";
            when "00" & x"020" => DATA <= x"003f";
            when "00" & x"021" => DATA <= x"0760";
            when "00" & x"022" => DATA <= x"003f";
            when "00" & x"023" => DATA <= x"0760";
            when "00" & x"024" => DATA <= x"003f";
            when "00" & x"025" => DATA <= x"0760";
            when "00" & x"026" => DATA <= x"003f";
            when "00" & x"027" => DATA <= x"0760";
            when "00" & x"028" => DATA <= x"003f";
            when "00" & x"029" => DATA <= x"0760";
            when "00" & x"02a" => DATA <= x"003f";
            when "00" & x"02b" => DATA <= x"0760";
            when "00" & x"02c" => DATA <= x"003f";
            when "00" & x"02d" => DATA <= x"0760";
            when "00" & x"02e" => DATA <= x"003f";
            when "00" & x"02f" => DATA <= x"0760";
            when "00" & x"030" => DATA <= x"003f";
            when "00" & x"031" => DATA <= x"0760";
            when "00" & x"032" => DATA <= x"003f";
            when "00" & x"033" => DATA <= x"25ae";
            when "00" & x"034" => DATA <= x"003f";
            when "00" & x"035" => DATA <= x"044c";
            when "00" & x"036" => DATA <= x"003f";
            when "00" & x"037" => DATA <= x"25ae";
            when "00" & x"038" => DATA <= x"003f";
            when "00" & x"039" => DATA <= x"25ae";
            when "00" & x"03a" => DATA <= x"003f";
            when "00" & x"03b" => DATA <= x"05fe";
            when "00" & x"03c" => DATA <= x"003f";
            when "00" & x"03d" => DATA <= x"25ae";
            when "00" & x"03e" => DATA <= x"003f";
            when "00" & x"03f" => DATA <= x"25ae";
            when "00" & x"040" => DATA <= x"003f";
            when "00" & x"041" => DATA <= x"0760";
            when "00" & x"042" => DATA <= x"003f";
            when "00" & x"043" => DATA <= x"0760";
            when "00" & x"044" => DATA <= x"003f";
            when "00" & x"045" => DATA <= x"0760";
            when "00" & x"046" => DATA <= x"003f";
            when "00" & x"047" => DATA <= x"0760";
            when "00" & x"048" => DATA <= x"003f";
            when "00" & x"049" => DATA <= x"0760";
            when "00" & x"04a" => DATA <= x"003f";
            when "00" & x"04b" => DATA <= x"0760";
            when "00" & x"04c" => DATA <= x"003f";
            when "00" & x"04d" => DATA <= x"0760";
            when "00" & x"04e" => DATA <= x"003f";
            when "00" & x"04f" => DATA <= x"0760";
            when "00" & x"050" => DATA <= x"003f";
            when "00" & x"051" => DATA <= x"0760";
            when "00" & x"052" => DATA <= x"003f";
            when "00" & x"053" => DATA <= x"0760";
            when "00" & x"054" => DATA <= x"003f";
            when "00" & x"055" => DATA <= x"0760";
            when "00" & x"056" => DATA <= x"003f";
            when "00" & x"057" => DATA <= x"0760";
            when "00" & x"058" => DATA <= x"003f";
            when "00" & x"059" => DATA <= x"08fc";
            when "00" & x"05a" => DATA <= x"003f";
            when "00" & x"05b" => DATA <= x"0760";
            when "00" & x"05c" => DATA <= x"003f";
            when "00" & x"05d" => DATA <= x"0760";
            when "00" & x"05e" => DATA <= x"003f";
            when "00" & x"05f" => DATA <= x"0760";
            when "00" & x"060" => DATA <= x"003f";
            when "00" & x"061" => DATA <= x"0760";
            when "00" & x"062" => DATA <= x"003f";
            when "00" & x"063" => DATA <= x"0760";
            when "00" & x"064" => DATA <= x"003f";
            when "00" & x"065" => DATA <= x"0760";
            when "00" & x"066" => DATA <= x"003f";
            when "00" & x"067" => DATA <= x"0760";
            when "00" & x"068" => DATA <= x"003f";
            when "00" & x"069" => DATA <= x"0760";
            when "00" & x"06a" => DATA <= x"003f";
            when "00" & x"06b" => DATA <= x"0760";
            when "00" & x"06c" => DATA <= x"003f";
            when "00" & x"06d" => DATA <= x"0760";
            when "00" & x"06e" => DATA <= x"003f";
            when "00" & x"06f" => DATA <= x"0760";
            when "00" & x"070" => DATA <= x"003f";
            when "00" & x"071" => DATA <= x"0760";
            when "00" & x"072" => DATA <= x"003f";
            when "00" & x"073" => DATA <= x"0760";
            when "00" & x"074" => DATA <= x"003f";
            when "00" & x"075" => DATA <= x"0760";
            when "00" & x"076" => DATA <= x"003f";
            when "00" & x"077" => DATA <= x"0760";
            when "00" & x"078" => DATA <= x"003f";
            when "00" & x"079" => DATA <= x"0760";
            when "00" & x"07a" => DATA <= x"003f";
            when "00" & x"07b" => DATA <= x"0760";
            when "00" & x"07c" => DATA <= x"003f";
            when "00" & x"07d" => DATA <= x"0760";
            when "00" & x"07e" => DATA <= x"003f";
            when "00" & x"07f" => DATA <= x"0760";
            when "00" & x"080" => DATA <= x"003f";
            when "00" & x"081" => DATA <= x"0776";
            when "00" & x"082" => DATA <= x"003f";
            when "00" & x"083" => DATA <= x"256c";
            when "00" & x"084" => DATA <= x"003f";
            when "00" & x"085" => DATA <= x"25ae";
            when "00" & x"086" => DATA <= x"003f";
            when "00" & x"087" => DATA <= x"25c6";
            when "00" & x"088" => DATA <= x"003f";
            when "00" & x"089" => DATA <= x"0a20";
            when "00" & x"08a" => DATA <= x"003f";
            when "00" & x"08b" => DATA <= x"0a30";
            when "00" & x"08c" => DATA <= x"003f";
            when "00" & x"08d" => DATA <= x"0ad2";
            when "00" & x"08e" => DATA <= x"003f";
            when "00" & x"08f" => DATA <= x"0be4";
            when "00" & x"090" => DATA <= x"003f";
            when "00" & x"091" => DATA <= x"0cca";
            when "00" & x"092" => DATA <= x"003f";
            when "00" & x"093" => DATA <= x"0d1a";
            when "00" & x"094" => DATA <= x"003f";
            when "00" & x"095" => DATA <= x"0d46";
            when "00" & x"096" => DATA <= x"003f";
            when "00" & x"097" => DATA <= x"0d5c";
            when "00" & x"098" => DATA <= x"003f";
            when "00" & x"099" => DATA <= x"0d7a";
            when "00" & x"09a" => DATA <= x"003f";
            when "00" & x"09b" => DATA <= x"0dbe";
            when "00" & x"09c" => DATA <= x"003f";
            when "00" & x"09d" => DATA <= x"0dec";
            when "00" & x"09e" => DATA <= x"003f";
            when "00" & x"09f" => DATA <= x"10d6";
            when "00" & x"0a0" => DATA <= x"003f";
            when "00" & x"0a1" => DATA <= x"25d8";
            when "00" & x"0a2" => DATA <= x"003f";
            when "00" & x"0a3" => DATA <= x"0776";
            when "00" & x"0a4" => DATA <= x"003f";
            when "00" & x"0a5" => DATA <= x"0776";
            when "00" & x"0a6" => DATA <= x"003f";
            when "00" & x"0a7" => DATA <= x"0776";
            when "00" & x"0a8" => DATA <= x"003f";
            when "00" & x"0a9" => DATA <= x"0776";
            when "00" & x"0aa" => DATA <= x"003f";
            when "00" & x"0ab" => DATA <= x"0776";
            when "00" & x"0ac" => DATA <= x"003f";
            when "00" & x"0ad" => DATA <= x"0776";
            when "00" & x"0ae" => DATA <= x"003f";
            when "00" & x"0af" => DATA <= x"0776";
            when "00" & x"0b0" => DATA <= x"003f";
            when "00" & x"0b1" => DATA <= x"25da";
            when "00" & x"0b2" => DATA <= x"003f";
            when "00" & x"0b3" => DATA <= x"0776";
            when "00" & x"0b4" => DATA <= x"003f";
            when "00" & x"0b5" => DATA <= x"0f0a";
            when "00" & x"0b6" => DATA <= x"003f";
            when "00" & x"0b7" => DATA <= x"0776";
            when "00" & x"0b8" => DATA <= x"003f";
            when "00" & x"0b9" => DATA <= x"0776";
            when "00" & x"0ba" => DATA <= x"003f";
            when "00" & x"0bb" => DATA <= x"0776";
            when "00" & x"0bc" => DATA <= x"003f";
            when "00" & x"0bd" => DATA <= x"25ea";
            when "00" & x"0be" => DATA <= x"003f";
            when "00" & x"0bf" => DATA <= x"0776";
            when "00" & x"0c0" => DATA <= x"003f";
            when "00" & x"0c1" => DATA <= x"0776";
            when "00" & x"0c2" => DATA <= x"003f";
            when "00" & x"0c3" => DATA <= x"0776";
            when "00" & x"0c4" => DATA <= x"003f";
            when "00" & x"0c5" => DATA <= x"0776";
            when "00" & x"0c6" => DATA <= x"003f";
            when "00" & x"0c7" => DATA <= x"0776";
            when "00" & x"0c8" => DATA <= x"003f";
            when "00" & x"0c9" => DATA <= x"0776";
            when "00" & x"0ca" => DATA <= x"003f";
            when "00" & x"0cb" => DATA <= x"0776";
            when "00" & x"0cc" => DATA <= x"003f";
            when "00" & x"0cd" => DATA <= x"0776";
            when "00" & x"0ce" => DATA <= x"003f";
            when "00" & x"0cf" => DATA <= x"0776";
            when "00" & x"0d0" => DATA <= x"003f";
            when "00" & x"0d1" => DATA <= x"0776";
            when "00" & x"0d2" => DATA <= x"003f";
            when "00" & x"0d3" => DATA <= x"0776";
            when "00" & x"0d4" => DATA <= x"003f";
            when "00" & x"0d5" => DATA <= x"0776";
            when "00" & x"0d6" => DATA <= x"003f";
            when "00" & x"0d7" => DATA <= x"0776";
            when "00" & x"0d8" => DATA <= x"0000";
            when "00" & x"0d9" => DATA <= x"0000";
            when "00" & x"0da" => DATA <= x"0000";
            when "00" & x"0db" => DATA <= x"0000";
            when "00" & x"0dc" => DATA <= x"0000";
            when "00" & x"0dd" => DATA <= x"0000";
            when "00" & x"0de" => DATA <= x"0000";
            when "00" & x"0df" => DATA <= x"0000";
            when "00" & x"0e0" => DATA <= x"0000";
            when "00" & x"0e1" => DATA <= x"0000";
            when "00" & x"0e2" => DATA <= x"003f";
            when "00" & x"0e3" => DATA <= x"2656";
            when "00" & x"0e4" => DATA <= x"003f";
            when "00" & x"0e5" => DATA <= x"265a";
            when "00" & x"0e6" => DATA <= x"003f";
            when "00" & x"0e7" => DATA <= x"265e";
            when "00" & x"0e8" => DATA <= x"003f";
            when "00" & x"0e9" => DATA <= x"2668";
            when "00" & x"0ea" => DATA <= x"0000";
            when "00" & x"0eb" => DATA <= x"0000";
            when "00" & x"0ec" => DATA <= x"0000";
            when "00" & x"0ed" => DATA <= x"0000";
            when "00" & x"0ee" => DATA <= x"0000";
            when "00" & x"0ef" => DATA <= x"0000";
            when "00" & x"0f0" => DATA <= x"0000";
            when "00" & x"0f1" => DATA <= x"0000";
            when "00" & x"0f2" => DATA <= x"0000";
            when "00" & x"0f3" => DATA <= x"0000";
            when "00" & x"0f4" => DATA <= x"0000";
            when "00" & x"0f5" => DATA <= x"0000";
            when "00" & x"0f6" => DATA <= x"0000";
            when "00" & x"0f7" => DATA <= x"0000";
            when "00" & x"0f8" => DATA <= x"0000";
            when "00" & x"0f9" => DATA <= x"0000";
            when "00" & x"0fa" => DATA <= x"0000";
            when "00" & x"0fb" => DATA <= x"0700";
            when "00" & x"0fc" => DATA <= x"0000";
            when "00" & x"0fd" => DATA <= x"0000";
            when "00" & x"0fe" => DATA <= x"0000";
            when "00" & x"0ff" => DATA <= x"0000";
            when "00" & x"100" => DATA <= x"207c";
            when "00" & x"101" => DATA <= x"0000";
            when "00" & x"102" => DATA <= x"0000";
            when "00" & x"103" => DATA <= x"227c";
            when "00" & x"104" => DATA <= x"003f";
            when "00" & x"105" => DATA <= x"0000";
            when "00" & x"106" => DATA <= x"303c";
            when "00" & x"107" => DATA <= x"003f";
            when "00" & x"108" => DATA <= x"20d9";
            when "00" & x"109" => DATA <= x"51c8";
            when "00" & x"10a" => DATA <= x"fffc";
            when "00" & x"10b" => DATA <= x"303c";
            when "00" & x"10c" => DATA <= x"00bf";
            when "00" & x"10d" => DATA <= x"20fc";
            when "00" & x"10e" => DATA <= x"003f";
            when "00" & x"10f" => DATA <= x"0760";
            when "00" & x"110" => DATA <= x"51c8";
            when "00" & x"111" => DATA <= x"fff8";
            when "00" & x"112" => DATA <= x"303c";
            when "00" & x"113" => DATA <= x"003f";
            when "00" & x"114" => DATA <= x"207c";
            when "00" & x"115" => DATA <= x"0000";
            when "00" & x"116" => DATA <= x"0400";
            when "00" & x"117" => DATA <= x"227c";
            when "00" & x"118" => DATA <= x"003f";
            when "00" & x"119" => DATA <= x"0100";
            when "00" & x"11a" => DATA <= x"20d9";
            when "00" & x"11b" => DATA <= x"51c8";
            when "00" & x"11c" => DATA <= x"fffc";
            when "00" & x"11d" => DATA <= x"203c";
            when "00" & x"11e" => DATA <= x"0001";
            when "00" & x"11f" => DATA <= x"fedf";
            when "00" & x"120" => DATA <= x"207c";
            when "00" & x"121" => DATA <= x"0000";
            when "00" & x"122" => DATA <= x"0500";
            when "00" & x"123" => DATA <= x"20fc";
            when "00" & x"124" => DATA <= x"0000";
            when "00" & x"125" => DATA <= x"0000";
            when "00" & x"126" => DATA <= x"51c8";
            when "00" & x"127" => DATA <= x"fff8";
            when "00" & x"128" => DATA <= x"6100";
            when "00" & x"129" => DATA <= x"0674";
            when "00" & x"12a" => DATA <= x"21c0";
            when "00" & x"12b" => DATA <= x"0508";
            when "00" & x"12c" => DATA <= x"2e40";
            when "00" & x"12d" => DATA <= x"0480";
            when "00" & x"12e" => DATA <= x"0000";
            when "00" & x"12f" => DATA <= x"0200";
            when "00" & x"130" => DATA <= x"2c40";
            when "00" & x"131" => DATA <= x"4e66";
            when "00" & x"132" => DATA <= x"0480";
            when "00" & x"133" => DATA <= x"0000";
            when "00" & x"134" => DATA <= x"0200";
            when "00" & x"135" => DATA <= x"23c0";
            when "00" & x"136" => DATA <= x"0000";
            when "00" & x"137" => DATA <= x"0500";
            when "00" & x"138" => DATA <= x"33fc";
            when "00" & x"139" => DATA <= x"0000";
            when "00" & x"13a" => DATA <= x"0000";
            when "00" & x"13b" => DATA <= x"0524";
            when "00" & x"13c" => DATA <= x"23fc";
            when "00" & x"13d" => DATA <= x"0000";
            when "00" & x"13e" => DATA <= x"0800";
            when "00" & x"13f" => DATA <= x"0000";
            when "00" & x"140" => DATA <= x"0504";
            when "00" & x"141" => DATA <= x"6100";
            when "00" & x"142" => DATA <= x"0502";
            when "00" & x"143" => DATA <= x"11c0";
            when "00" & x"144" => DATA <= x"0532";
            when "00" & x"145" => DATA <= x"6100";
            when "00" & x"146" => DATA <= x"0578";
            when "00" & x"147" => DATA <= x"11c0";
            when "00" & x"148" => DATA <= x"0533";
            when "00" & x"149" => DATA <= x"6100";
            when "00" & x"14a" => DATA <= x"0592";
            when "00" & x"14b" => DATA <= x"11c0";
            when "00" & x"14c" => DATA <= x"0534";
            when "00" & x"14d" => DATA <= x"11fc";
            when "00" & x"14e" => DATA <= x"0000";
            when "00" & x"14f" => DATA <= x"0535";
            when "00" & x"150" => DATA <= x"027c";
            when "00" & x"151" => DATA <= x"dfff";
            when "00" & x"152" => DATA <= x"203c";
            when "00" & x"153" => DATA <= x"003f";
            when "00" & x"154" => DATA <= x"27e2";
            when "00" & x"155" => DATA <= x"6100";
            when "00" & x"156" => DATA <= x"0752";
            when "00" & x"157" => DATA <= x"1038";
            when "00" & x"158" => DATA <= x"0532";
            when "00" & x"159" => DATA <= x"b07c";
            when "00" & x"15a" => DATA <= x"0009";
            when "00" & x"15b" => DATA <= x"6500";
            when "00" & x"15c" => DATA <= x"0004";
            when "00" & x"15d" => DATA <= x"7000";
            when "00" & x"15e" => DATA <= x"0c38";
            when "00" & x"15f" => DATA <= x"00ff";
            when "00" & x"160" => DATA <= x"0532";
            when "00" & x"161" => DATA <= x"6700";
            when "00" & x"162" => DATA <= x"001e";
            when "00" & x"163" => DATA <= x"203c";
            when "00" & x"164" => DATA <= x"003f";
            when "00" & x"165" => DATA <= x"2800";
            when "00" & x"166" => DATA <= x"d038";
            when "00" & x"167" => DATA <= x"0532";
            when "00" & x"168" => DATA <= x"d038";
            when "00" & x"169" => DATA <= x"0532";
            when "00" & x"16a" => DATA <= x"d038";
            when "00" & x"16b" => DATA <= x"0532";
            when "00" & x"16c" => DATA <= x"7203";
            when "00" & x"16d" => DATA <= x"6100";
            when "00" & x"16e" => DATA <= x"1092";
            when "00" & x"16f" => DATA <= x"6000";
            when "00" & x"170" => DATA <= x"000a";
            when "00" & x"171" => DATA <= x"103c";
            when "00" & x"172" => DATA <= x"004b";
            when "00" & x"173" => DATA <= x"6100";
            when "00" & x"174" => DATA <= x"06fe";
            when "00" & x"175" => DATA <= x"203c";
            when "00" & x"176" => DATA <= x"003f";
            when "00" & x"177" => DATA <= x"27ed";
            when "00" & x"178" => DATA <= x"6100";
            when "00" & x"179" => DATA <= x"070c";
            when "00" & x"17a" => DATA <= x"2038";
            when "00" & x"17b" => DATA <= x"0508";
            when "00" & x"17c" => DATA <= x"ea88";
            when "00" & x"17d" => DATA <= x"ea88";
            when "00" & x"17e" => DATA <= x"223c";
            when "00" & x"17f" => DATA <= x"0000";
            when "00" & x"180" => DATA <= x"0600";
            when "00" & x"181" => DATA <= x"243c";
            when "00" & x"182" => DATA <= x"0000";
            when "00" & x"183" => DATA <= x"00ff";
            when "00" & x"184" => DATA <= x"6100";
            when "00" & x"185" => DATA <= x"1484";
            when "00" & x"186" => DATA <= x"203c";
            when "00" & x"187" => DATA <= x"0000";
            when "00" & x"188" => DATA <= x"0600";
            when "00" & x"189" => DATA <= x"6100";
            when "00" & x"18a" => DATA <= x"06ea";
            when "00" & x"18b" => DATA <= x"203c";
            when "00" & x"18c" => DATA <= x"003f";
            when "00" & x"18d" => DATA <= x"281b";
            when "00" & x"18e" => DATA <= x"7207";
            when "00" & x"18f" => DATA <= x"6100";
            when "00" & x"190" => DATA <= x"104e";
            when "00" & x"191" => DATA <= x"7227";
            when "00" & x"192" => DATA <= x"6100";
            when "00" & x"193" => DATA <= x"0e2a";
            when "00" & x"194" => DATA <= x"6100";
            when "00" & x"195" => DATA <= x"00a6";
            when "00" & x"196" => DATA <= x"2f00";
            when "00" & x"197" => DATA <= x"7001";
            when "00" & x"198" => DATA <= x"223c";
            when "00" & x"199" => DATA <= x"0000";
            when "00" & x"19a" => DATA <= x"0528";
            when "00" & x"19b" => DATA <= x"6100";
            when "00" & x"19c" => DATA <= x"08ac";
            when "00" & x"19d" => DATA <= x"11fc";
            when "00" & x"19e" => DATA <= x"0000";
            when "00" & x"19f" => DATA <= x"052d";
            when "00" & x"1a0" => DATA <= x"11fc";
            when "00" & x"1a1" => DATA <= x"0000";
            when "00" & x"1a2" => DATA <= x"052e";
            when "00" & x"1a3" => DATA <= x"11fc";
            when "00" & x"1a4" => DATA <= x"0000";
            when "00" & x"1a5" => DATA <= x"052f";
            when "00" & x"1a6" => DATA <= x"11fc";
            when "00" & x"1a7" => DATA <= x"0000";
            when "00" & x"1a8" => DATA <= x"0530";
            when "00" & x"1a9" => DATA <= x"11fc";
            when "00" & x"1aa" => DATA <= x"0000";
            when "00" & x"1ab" => DATA <= x"0531";
            when "00" & x"1ac" => DATA <= x"201f";
            when "00" & x"1ad" => DATA <= x"b03c";
            when "00" & x"1ae" => DATA <= x"0080";
            when "00" & x"1af" => DATA <= x"103c";
            when "00" & x"1b0" => DATA <= x"002a";
            when "00" & x"1b1" => DATA <= x"6100";
            when "00" & x"1b2" => DATA <= x"0682";
            when "00" & x"1b3" => DATA <= x"203c";
            when "00" & x"1b4" => DATA <= x"0000";
            when "00" & x"1b5" => DATA <= x"0600";
            when "00" & x"1b6" => DATA <= x"223c";
            when "00" & x"1b7" => DATA <= x"0000";
            when "00" & x"1b8" => DATA <= x"00ff";
            when "00" & x"1b9" => DATA <= x"143c";
            when "00" & x"1ba" => DATA <= x"0020";
            when "00" & x"1bb" => DATA <= x"163c";
            when "00" & x"1bc" => DATA <= x"00ff";
            when "00" & x"1bd" => DATA <= x"207c";
            when "00" & x"1be" => DATA <= x"0000";
            when "00" & x"1bf" => DATA <= x"007d";
            when "00" & x"1c0" => DATA <= x"4e4c";
            when "00" & x"1c1" => DATA <= x"6500";
            when "00" & x"1c2" => DATA <= x"0012";
            when "00" & x"1c3" => DATA <= x"203c";
            when "00" & x"1c4" => DATA <= x"0000";
            when "00" & x"1c5" => DATA <= x"0600";
            when "00" & x"1c6" => DATA <= x"207c";
            when "00" & x"1c7" => DATA <= x"0000";
            when "00" & x"1c8" => DATA <= x"0005";
            when "00" & x"1c9" => DATA <= x"4e4c";
            when "00" & x"1ca" => DATA <= x"60c8";
            when "00" & x"1cb" => DATA <= x"707e";
            when "00" & x"1cc" => DATA <= x"6100";
            when "00" & x"1cd" => DATA <= x"0738";
            when "00" & x"1ce" => DATA <= x"203c";
            when "00" & x"1cf" => DATA <= x"003f";
            when "00" & x"1d0" => DATA <= x"2d78";
            when "00" & x"1d1" => DATA <= x"207c";
            when "00" & x"1d2" => DATA <= x"0000";
            when "00" & x"1d3" => DATA <= x"002b";
            when "00" & x"1d4" => DATA <= x"4e4c";
            when "00" & x"1d5" => DATA <= x"60b2";
            when "00" & x"1d6" => DATA <= x"0839";
            when "00" & x"1d7" => DATA <= x"0007";
            when "00" & x"1d8" => DATA <= x"fffe";
            when "00" & x"1d9" => DATA <= x"0000";
            when "00" & x"1da" => DATA <= x"6600";
            when "00" & x"1db" => DATA <= x"0012";
            when "00" & x"1dc" => DATA <= x"0839";
            when "00" & x"1dd" => DATA <= x"0007";
            when "00" & x"1de" => DATA <= x"fffe";
            when "00" & x"1df" => DATA <= x"0006";
            when "00" & x"1e0" => DATA <= x"67ea";
            when "00" & x"1e1" => DATA <= x"6100";
            when "00" & x"1e2" => DATA <= x"00f0";
            when "00" & x"1e3" => DATA <= x"60e4";
            when "00" & x"1e4" => DATA <= x"1039";
            when "00" & x"1e5" => DATA <= x"fffe";
            when "00" & x"1e6" => DATA <= x"0001";
            when "00" & x"1e7" => DATA <= x"4e75";
            when "00" & x"1e8" => DATA <= x"0839";
            when "00" & x"1e9" => DATA <= x"0007";
            when "00" & x"1ea" => DATA <= x"fffe";
            when "00" & x"1eb" => DATA <= x"0002";
            when "00" & x"1ec" => DATA <= x"67f6";
            when "00" & x"1ed" => DATA <= x"1039";
            when "00" & x"1ee" => DATA <= x"fffe";
            when "00" & x"1ef" => DATA <= x"0003";
            when "00" & x"1f0" => DATA <= x"4e75";
            when "00" & x"1f1" => DATA <= x"0839";
            when "00" & x"1f2" => DATA <= x"0006";
            when "00" & x"1f3" => DATA <= x"fffe";
            when "00" & x"1f4" => DATA <= x"0002";
            when "00" & x"1f5" => DATA <= x"67f6";
            when "00" & x"1f6" => DATA <= x"13c0";
            when "00" & x"1f7" => DATA <= x"fffe";
            when "00" & x"1f8" => DATA <= x"0003";
            when "00" & x"1f9" => DATA <= x"4e75";
            when "00" & x"1fa" => DATA <= x"0839";
            when "00" & x"1fb" => DATA <= x"0007";
            when "00" & x"1fc" => DATA <= x"fffe";
            when "00" & x"1fd" => DATA <= x"0006";
            when "00" & x"1fe" => DATA <= x"67f6";
            when "00" & x"1ff" => DATA <= x"1039";
            when "00" & x"200" => DATA <= x"fffe";
            when "00" & x"201" => DATA <= x"0007";
            when "00" & x"202" => DATA <= x"4e75";
            when "00" & x"203" => DATA <= x"4280";
            when "00" & x"204" => DATA <= x"61c6";
            when "00" & x"205" => DATA <= x"e198";
            when "00" & x"206" => DATA <= x"61c2";
            when "00" & x"207" => DATA <= x"e198";
            when "00" & x"208" => DATA <= x"61be";
            when "00" & x"209" => DATA <= x"e198";
            when "00" & x"20a" => DATA <= x"60ba";
            when "00" & x"20b" => DATA <= x"e198";
            when "00" & x"20c" => DATA <= x"61c8";
            when "00" & x"20d" => DATA <= x"e198";
            when "00" & x"20e" => DATA <= x"61c4";
            when "00" & x"20f" => DATA <= x"e198";
            when "00" & x"210" => DATA <= x"61c0";
            when "00" & x"211" => DATA <= x"e198";
            when "00" & x"212" => DATA <= x"60bc";
            when "00" & x"213" => DATA <= x"4280";
            when "00" & x"214" => DATA <= x"61ca";
            when "00" & x"215" => DATA <= x"e198";
            when "00" & x"216" => DATA <= x"61c6";
            when "00" & x"217" => DATA <= x"e198";
            when "00" & x"218" => DATA <= x"61c2";
            when "00" & x"219" => DATA <= x"e198";
            when "00" & x"21a" => DATA <= x"60be";
            when "00" & x"21b" => DATA <= x"0839";
            when "00" & x"21c" => DATA <= x"0006";
            when "00" & x"21d" => DATA <= x"fffe";
            when "00" & x"21e" => DATA <= x"0002";
            when "00" & x"21f" => DATA <= x"67f6";
            when "00" & x"220" => DATA <= x"101e";
            when "00" & x"221" => DATA <= x"619e";
            when "00" & x"222" => DATA <= x"b03c";
            when "00" & x"223" => DATA <= x"000d";
            when "00" & x"224" => DATA <= x"66ec";
            when "00" & x"225" => DATA <= x"4e75";
            when "00" & x"226" => DATA <= x"0839";
            when "00" & x"227" => DATA <= x"0007";
            when "00" & x"228" => DATA <= x"fffe";
            when "00" & x"229" => DATA <= x"0006";
            when "00" & x"22a" => DATA <= x"6600";
            when "00" & x"22b" => DATA <= x"005e";
            when "00" & x"22c" => DATA <= x"0839";
            when "00" & x"22d" => DATA <= x"0007";
            when "00" & x"22e" => DATA <= x"fffe";
            when "00" & x"22f" => DATA <= x"0000";
            when "00" & x"230" => DATA <= x"6600";
            when "00" & x"231" => DATA <= x"0010";
            when "00" & x"232" => DATA <= x"2f0e";
            when "00" & x"233" => DATA <= x"2c79";
            when "00" & x"234" => DATA <= x"0000";
            when "00" & x"235" => DATA <= x"0408";
            when "00" & x"236" => DATA <= x"4e96";
            when "00" & x"237" => DATA <= x"2c5f";
            when "00" & x"238" => DATA <= x"4e73";
            when "00" & x"239" => DATA <= x"2f00";
            when "00" & x"23a" => DATA <= x"1039";
            when "00" & x"23b" => DATA <= x"fffe";
            when "00" & x"23c" => DATA <= x"0001";
            when "00" & x"23d" => DATA <= x"6b00";
            when "00" & x"23e" => DATA <= x"0028";
            when "00" & x"23f" => DATA <= x"2f01";
            when "00" & x"240" => DATA <= x"4280";
            when "00" & x"241" => DATA <= x"6100";
            when "00" & x"242" => DATA <= x"ff28";
            when "00" & x"243" => DATA <= x"e158";
            when "00" & x"244" => DATA <= x"6100";
            when "00" & x"245" => DATA <= x"ff22";
            when "00" & x"246" => DATA <= x"3200";
            when "00" & x"247" => DATA <= x"6100";
            when "00" & x"248" => DATA <= x"ff1c";
            when "00" & x"249" => DATA <= x"2f0e";
            when "00" & x"24a" => DATA <= x"2c79";
            when "00" & x"24b" => DATA <= x"0000";
            when "00" & x"24c" => DATA <= x"0440";
            when "00" & x"24d" => DATA <= x"4e96";
            when "00" & x"24e" => DATA <= x"2c5f";
            when "00" & x"24f" => DATA <= x"221f";
            when "00" & x"250" => DATA <= x"201f";
            when "00" & x"251" => DATA <= x"4e73";
            when "00" & x"252" => DATA <= x"2f0e";
            when "00" & x"253" => DATA <= x"2c79";
            when "00" & x"254" => DATA <= x"0000";
            when "00" & x"255" => DATA <= x"04cc";
            when "00" & x"256" => DATA <= x"4e96";
            when "00" & x"257" => DATA <= x"2c5f";
            when "00" & x"258" => DATA <= x"201f";
            when "00" & x"259" => DATA <= x"4e73";
            when "00" & x"25a" => DATA <= x"1039";
            when "00" & x"25b" => DATA <= x"fffe";
            when "00" & x"25c" => DATA <= x"0007";
            when "00" & x"25d" => DATA <= x"6a00";
            when "00" & x"25e" => DATA <= x"003c";
            when "00" & x"25f" => DATA <= x"2f00";
            when "00" & x"260" => DATA <= x"2f0e";
            when "00" & x"261" => DATA <= x"2c7c";
            when "00" & x"262" => DATA <= x"0000";
            when "00" & x"263" => DATA <= x"0700";
            when "00" & x"264" => DATA <= x"6100";
            when "00" & x"265" => DATA <= x"ff06";
            when "00" & x"266" => DATA <= x"4280";
            when "00" & x"267" => DATA <= x"6100";
            when "00" & x"268" => DATA <= x"ff00";
            when "00" & x"269" => DATA <= x"2cc0";
            when "00" & x"26a" => DATA <= x"6100";
            when "00" & x"26b" => DATA <= x"fefa";
            when "00" & x"26c" => DATA <= x"1cc0";
            when "00" & x"26d" => DATA <= x"66f8";
            when "00" & x"26e" => DATA <= x"2c5f";
            when "00" & x"26f" => DATA <= x"203c";
            when "00" & x"270" => DATA <= x"0000";
            when "00" & x"271" => DATA <= x"0700";
            when "00" & x"272" => DATA <= x"21c0";
            when "00" & x"273" => DATA <= x"0514";
            when "00" & x"274" => DATA <= x"21fc";
            when "00" & x"275" => DATA <= x"ffff";
            when "00" & x"276" => DATA <= x"6502";
            when "00" & x"277" => DATA <= x"0510";
            when "00" & x"278" => DATA <= x"6100";
            when "00" & x"279" => DATA <= x"0c2e";
            when "00" & x"27a" => DATA <= x"201f";
            when "00" & x"27b" => DATA <= x"4e73";
            when "00" & x"27c" => DATA <= x"2f08";
            when "00" & x"27d" => DATA <= x"2f00";
            when "00" & x"27e" => DATA <= x"0280";
            when "00" & x"27f" => DATA <= x"0000";
            when "00" & x"280" => DATA <= x"00ff";
            when "00" & x"281" => DATA <= x"e588";
            when "00" & x"282" => DATA <= x"41f9";
            when "00" & x"283" => DATA <= x"003f";
            when "00" & x"284" => DATA <= x"0606";
            when "00" & x"285" => DATA <= x"d1c0";
            when "00" & x"286" => DATA <= x"21c8";
            when "00" & x"287" => DATA <= x"0074";
            when "00" & x"288" => DATA <= x"6100";
            when "00" & x"289" => DATA <= x"fee2";
            when "00" & x"28a" => DATA <= x"2017";
            when "00" & x"28b" => DATA <= x"b03c";
            when "00" & x"28c" => DATA <= x"0005";
            when "00" & x"28d" => DATA <= x"6700";
            when "00" & x"28e" => DATA <= x"005c";
            when "00" & x"28f" => DATA <= x"6100";
            when "00" & x"290" => DATA <= x"ff06";
            when "00" & x"291" => DATA <= x"23c0";
            when "00" & x"292" => DATA <= x"0000";
            when "00" & x"293" => DATA <= x"0520";
            when "00" & x"294" => DATA <= x"1039";
            when "00" & x"295" => DATA <= x"fffe";
            when "00" & x"296" => DATA <= x"0005";
            when "00" & x"297" => DATA <= x"1039";
            when "00" & x"298" => DATA <= x"fffe";
            when "00" & x"299" => DATA <= x"0005";
            when "00" & x"29a" => DATA <= x"6100";
            when "00" & x"29b" => DATA <= x"febe";
            when "00" & x"29c" => DATA <= x"2017";
            when "00" & x"29d" => DATA <= x"b03c";
            when "00" & x"29e" => DATA <= x"0006";
            when "00" & x"29f" => DATA <= x"6500";
            when "00" & x"2a0" => DATA <= x"0038";
            when "00" & x"2a1" => DATA <= x"6600";
            when "00" & x"2a2" => DATA <= x"003a";
            when "00" & x"2a3" => DATA <= x"2f0e";
            when "00" & x"2a4" => DATA <= x"2c78";
            when "00" & x"2a5" => DATA <= x"0520";
            when "00" & x"2a6" => DATA <= x"203c";
            when "00" & x"2a7" => DATA <= x"0000";
            when "00" & x"2a8" => DATA <= x"00ff";
            when "00" & x"2a9" => DATA <= x"0839";
            when "00" & x"2aa" => DATA <= x"0007";
            when "00" & x"2ab" => DATA <= x"fffe";
            when "00" & x"2ac" => DATA <= x"0004";
            when "00" & x"2ad" => DATA <= x"67f6";
            when "00" & x"2ae" => DATA <= x"13de";
            when "00" & x"2af" => DATA <= x"fffe";
            when "00" & x"2b0" => DATA <= x"0005";
            when "00" & x"2b1" => DATA <= x"51c8";
            when "00" & x"2b2" => DATA <= x"ffee";
            when "00" & x"2b3" => DATA <= x"0839";
            when "00" & x"2b4" => DATA <= x"0007";
            when "00" & x"2b5" => DATA <= x"fffe";
            when "00" & x"2b6" => DATA <= x"0004";
            when "00" & x"2b7" => DATA <= x"67f6";
            when "00" & x"2b8" => DATA <= x"13e6";
            when "00" & x"2b9" => DATA <= x"fffe";
            when "00" & x"2ba" => DATA <= x"0005";
            when "00" & x"2bb" => DATA <= x"2c5f";
            when "00" & x"2bc" => DATA <= x"201f";
            when "00" & x"2bd" => DATA <= x"205f";
            when "00" & x"2be" => DATA <= x"4e73";
            when "00" & x"2bf" => DATA <= x"2f0e";
            when "00" & x"2c0" => DATA <= x"2c78";
            when "00" & x"2c1" => DATA <= x"0520";
            when "00" & x"2c2" => DATA <= x"203c";
            when "00" & x"2c3" => DATA <= x"0000";
            when "00" & x"2c4" => DATA <= x"00ff";
            when "00" & x"2c5" => DATA <= x"0839";
            when "00" & x"2c6" => DATA <= x"0007";
            when "00" & x"2c7" => DATA <= x"fffe";
            when "00" & x"2c8" => DATA <= x"0004";
            when "00" & x"2c9" => DATA <= x"67f6";
            when "00" & x"2ca" => DATA <= x"1cf9";
            when "00" & x"2cb" => DATA <= x"fffe";
            when "00" & x"2cc" => DATA <= x"0005";
            when "00" & x"2cd" => DATA <= x"51c8";
            when "00" & x"2ce" => DATA <= x"ffee";
            when "00" & x"2cf" => DATA <= x"2c5f";
            when "00" & x"2d0" => DATA <= x"60d6";
            when "00" & x"2d1" => DATA <= x"2f0e";
            when "00" & x"2d2" => DATA <= x"2c78";
            when "00" & x"2d3" => DATA <= x"0520";
            when "00" & x"2d4" => DATA <= x"13de";
            when "00" & x"2d5" => DATA <= x"fffe";
            when "00" & x"2d6" => DATA <= x"0005";
            when "00" & x"2d7" => DATA <= x"21ce";
            when "00" & x"2d8" => DATA <= x"0520";
            when "00" & x"2d9" => DATA <= x"2c5f";
            when "00" & x"2da" => DATA <= x"4e73";
            when "00" & x"2db" => DATA <= x"2f0e";
            when "00" & x"2dc" => DATA <= x"2c78";
            when "00" & x"2dd" => DATA <= x"0520";
            when "00" & x"2de" => DATA <= x"1cf9";
            when "00" & x"2df" => DATA <= x"fffe";
            when "00" & x"2e0" => DATA <= x"0005";
            when "00" & x"2e1" => DATA <= x"21ce";
            when "00" & x"2e2" => DATA <= x"0520";
            when "00" & x"2e3" => DATA <= x"2c5f";
            when "00" & x"2e4" => DATA <= x"4e73";
            when "00" & x"2e5" => DATA <= x"2f0e";
            when "00" & x"2e6" => DATA <= x"2c78";
            when "00" & x"2e7" => DATA <= x"0520";
            when "00" & x"2e8" => DATA <= x"13de";
            when "00" & x"2e9" => DATA <= x"fffe";
            when "00" & x"2ea" => DATA <= x"0005";
            when "00" & x"2eb" => DATA <= x"13de";
            when "00" & x"2ec" => DATA <= x"fffe";
            when "00" & x"2ed" => DATA <= x"0005";
            when "00" & x"2ee" => DATA <= x"21ce";
            when "00" & x"2ef" => DATA <= x"0520";
            when "00" & x"2f0" => DATA <= x"2c5f";
            when "00" & x"2f1" => DATA <= x"4e73";
            when "00" & x"2f2" => DATA <= x"2f0e";
            when "00" & x"2f3" => DATA <= x"2c78";
            when "00" & x"2f4" => DATA <= x"0520";
            when "00" & x"2f5" => DATA <= x"1cf9";
            when "00" & x"2f6" => DATA <= x"fffe";
            when "00" & x"2f7" => DATA <= x"0005";
            when "00" & x"2f8" => DATA <= x"1cf9";
            when "00" & x"2f9" => DATA <= x"fffe";
            when "00" & x"2fa" => DATA <= x"0005";
            when "00" & x"2fb" => DATA <= x"21ce";
            when "00" & x"2fc" => DATA <= x"0520";
            when "00" & x"2fd" => DATA <= x"2c5f";
            when "00" & x"2fe" => DATA <= x"4e73";
            when "00" & x"2ff" => DATA <= x"13c0";
            when "00" & x"300" => DATA <= x"fffe";
            when "00" & x"301" => DATA <= x"0005";
            when "00" & x"302" => DATA <= x"4e73";
            when "00" & x"303" => DATA <= x"003f";
            when "00" & x"304" => DATA <= x"05a2";
            when "00" & x"305" => DATA <= x"003f";
            when "00" & x"306" => DATA <= x"05b6";
            when "00" & x"307" => DATA <= x"003f";
            when "00" & x"308" => DATA <= x"05ca";
            when "00" & x"309" => DATA <= x"003f";
            when "00" & x"30a" => DATA <= x"05e4";
            when "00" & x"30b" => DATA <= x"003f";
            when "00" & x"30c" => DATA <= x"05fe";
            when "00" & x"30d" => DATA <= x"003f";
            when "00" & x"30e" => DATA <= x"05fe";
            when "00" & x"30f" => DATA <= x"003f";
            when "00" & x"310" => DATA <= x"05fe";
            when "00" & x"311" => DATA <= x"003f";
            when "00" & x"312" => DATA <= x"05fe";
            when "00" & x"313" => DATA <= x"203c";
            when "00" & x"314" => DATA <= x"003f";
            when "00" & x"315" => DATA <= x"2c49";
            when "00" & x"316" => DATA <= x"6100";
            when "00" & x"317" => DATA <= x"03d0";
            when "00" & x"318" => DATA <= x"31df";
            when "00" & x"319" => DATA <= x"0544";
            when "00" & x"31a" => DATA <= x"21df";
            when "00" & x"31b" => DATA <= x"0540";
            when "00" & x"31c" => DATA <= x"31df";
            when "00" & x"31d" => DATA <= x"053e";
            when "00" & x"31e" => DATA <= x"31df";
            when "00" & x"31f" => DATA <= x"053c";
            when "00" & x"320" => DATA <= x"21d7";
            when "00" & x"321" => DATA <= x"0538";
            when "00" & x"322" => DATA <= x"223c";
            when "00" & x"323" => DATA <= x"0000";
            when "00" & x"324" => DATA <= x"0600";
            when "00" & x"325" => DATA <= x"143c";
            when "00" & x"326" => DATA <= x"00ff";
            when "00" & x"327" => DATA <= x"7000";
            when "00" & x"328" => DATA <= x"2038";
            when "00" & x"329" => DATA <= x"0538";
            when "00" & x"32a" => DATA <= x"6100";
            when "00" & x"32b" => DATA <= x"1090";
            when "00" & x"32c" => DATA <= x"6100";
            when "00" & x"32d" => DATA <= x"03a4";
            when "00" & x"32e" => DATA <= x"6100";
            when "00" & x"32f" => DATA <= x"03b4";
            when "00" & x"330" => DATA <= x"203c";
            when "00" & x"331" => DATA <= x"003f";
            when "00" & x"332" => DATA <= x"2c79";
            when "00" & x"333" => DATA <= x"6100";
            when "00" & x"334" => DATA <= x"0396";
            when "00" & x"335" => DATA <= x"223c";
            when "00" & x"336" => DATA <= x"0000";
            when "00" & x"337" => DATA <= x"0600";
            when "00" & x"338" => DATA <= x"143c";
            when "00" & x"339" => DATA <= x"00ff";
            when "00" & x"33a" => DATA <= x"7000";
            when "00" & x"33b" => DATA <= x"3038";
            when "00" & x"33c" => DATA <= x"0544";
            when "00" & x"33d" => DATA <= x"6100";
            when "00" & x"33e" => DATA <= x"1030";
            when "00" & x"33f" => DATA <= x"6100";
            when "00" & x"340" => DATA <= x"037e";
            when "00" & x"341" => DATA <= x"6100";
            when "00" & x"342" => DATA <= x"038e";
            when "00" & x"343" => DATA <= x"203c";
            when "00" & x"344" => DATA <= x"003f";
            when "00" & x"345" => DATA <= x"2c90";
            when "00" & x"346" => DATA <= x"6100";
            when "00" & x"347" => DATA <= x"0370";
            when "00" & x"348" => DATA <= x"223c";
            when "00" & x"349" => DATA <= x"0000";
            when "00" & x"34a" => DATA <= x"0600";
            when "00" & x"34b" => DATA <= x"143c";
            when "00" & x"34c" => DATA <= x"00ff";
            when "00" & x"34d" => DATA <= x"7000";
            when "00" & x"34e" => DATA <= x"2038";
            when "00" & x"34f" => DATA <= x"0540";
            when "00" & x"350" => DATA <= x"6100";
            when "00" & x"351" => DATA <= x"1044";
            when "00" & x"352" => DATA <= x"6100";
            when "00" & x"353" => DATA <= x"0358";
            when "00" & x"354" => DATA <= x"6100";
            when "00" & x"355" => DATA <= x"0368";
            when "00" & x"356" => DATA <= x"203c";
            when "00" & x"357" => DATA <= x"003f";
            when "00" & x"358" => DATA <= x"2ca7";
            when "00" & x"359" => DATA <= x"6100";
            when "00" & x"35a" => DATA <= x"034a";
            when "00" & x"35b" => DATA <= x"223c";
            when "00" & x"35c" => DATA <= x"0000";
            when "00" & x"35d" => DATA <= x"0600";
            when "00" & x"35e" => DATA <= x"143c";
            when "00" & x"35f" => DATA <= x"00ff";
            when "00" & x"360" => DATA <= x"7000";
            when "00" & x"361" => DATA <= x"3038";
            when "00" & x"362" => DATA <= x"053e";
            when "00" & x"363" => DATA <= x"6100";
            when "00" & x"364" => DATA <= x"0fe4";
            when "00" & x"365" => DATA <= x"6100";
            when "00" & x"366" => DATA <= x"0332";
            when "00" & x"367" => DATA <= x"103c";
            when "00" & x"368" => DATA <= x"0020";
            when "00" & x"369" => DATA <= x"6100";
            when "00" & x"36a" => DATA <= x"0312";
            when "00" & x"36b" => DATA <= x"103c";
            when "00" & x"36c" => DATA <= x"005b";
            when "00" & x"36d" => DATA <= x"6100";
            when "00" & x"36e" => DATA <= x"030a";
            when "00" & x"36f" => DATA <= x"303c";
            when "00" & x"370" => DATA <= x"053e";
            when "00" & x"371" => DATA <= x"223c";
            when "00" & x"372" => DATA <= x"0000";
            when "00" & x"373" => DATA <= x"0600";
            when "00" & x"374" => DATA <= x"6100";
            when "00" & x"375" => DATA <= x"1422";
            when "00" & x"376" => DATA <= x"2001";
            when "00" & x"377" => DATA <= x"6100";
            when "00" & x"378" => DATA <= x"030e";
            when "00" & x"379" => DATA <= x"103c";
            when "00" & x"37a" => DATA <= x"005d";
            when "00" & x"37b" => DATA <= x"6100";
            when "00" & x"37c" => DATA <= x"02ee";
            when "00" & x"37d" => DATA <= x"6100";
            when "00" & x"37e" => DATA <= x"0316";
            when "00" & x"37f" => DATA <= x"203c";
            when "00" & x"380" => DATA <= x"003f";
            when "00" & x"381" => DATA <= x"2cbe";
            when "00" & x"382" => DATA <= x"6100";
            when "00" & x"383" => DATA <= x"02f8";
            when "00" & x"384" => DATA <= x"223c";
            when "00" & x"385" => DATA <= x"0000";
            when "00" & x"386" => DATA <= x"0600";
            when "00" & x"387" => DATA <= x"143c";
            when "00" & x"388" => DATA <= x"00ff";
            when "00" & x"389" => DATA <= x"7000";
            when "00" & x"38a" => DATA <= x"3038";
            when "00" & x"38b" => DATA <= x"053c";
            when "00" & x"38c" => DATA <= x"6100";
            when "00" & x"38d" => DATA <= x"120e";
            when "00" & x"38e" => DATA <= x"6100";
            when "00" & x"38f" => DATA <= x"02e0";
            when "00" & x"390" => DATA <= x"6100";
            when "00" & x"391" => DATA <= x"02f0";
            when "00" & x"392" => DATA <= x"60fe";
            when "00" & x"393" => DATA <= x"6100";
            when "00" & x"394" => DATA <= x"02f8";
            when "00" & x"395" => DATA <= x"6000";
            when "00" & x"396" => DATA <= x"fc32";
            when "00" & x"397" => DATA <= x"203c";
            when "00" & x"398" => DATA <= x"003f";
            when "00" & x"399" => DATA <= x"2c5a";
            when "00" & x"39a" => DATA <= x"6100";
            when "00" & x"39b" => DATA <= x"02c8";
            when "00" & x"39c" => DATA <= x"6000";
            when "00" & x"39d" => DATA <= x"fef6";
            when "00" & x"39e" => DATA <= x"2f00";
            when "00" & x"39f" => DATA <= x"203c";
            when "00" & x"3a0" => DATA <= x"003f";
            when "00" & x"3a1" => DATA <= x"2d00";
            when "00" & x"3a2" => DATA <= x"6000";
            when "00" & x"3a3" => DATA <= x"0022";
            when "00" & x"3a4" => DATA <= x"2f00";
            when "00" & x"3a5" => DATA <= x"203c";
            when "00" & x"3a6" => DATA <= x"003f";
            when "00" & x"3a7" => DATA <= x"2d30";
            when "00" & x"3a8" => DATA <= x"6000";
            when "00" & x"3a9" => DATA <= x"0016";
            when "00" & x"3aa" => DATA <= x"2f00";
            when "00" & x"3ab" => DATA <= x"203c";
            when "00" & x"3ac" => DATA <= x"003f";
            when "00" & x"3ad" => DATA <= x"2d4c";
            when "00" & x"3ae" => DATA <= x"6000";
            when "00" & x"3af" => DATA <= x"000a";
            when "00" & x"3b0" => DATA <= x"2f00";
            when "00" & x"3b1" => DATA <= x"203c";
            when "00" & x"3b2" => DATA <= x"003f";
            when "00" & x"3b3" => DATA <= x"2dbc";
            when "00" & x"3b4" => DATA <= x"21ef";
            when "00" & x"3b5" => DATA <= x"0006";
            when "00" & x"3b6" => DATA <= x"0510";
            when "00" & x"3b7" => DATA <= x"6100";
            when "00" & x"3b8" => DATA <= x"09b0";
            when "00" & x"3b9" => DATA <= x"201f";
            when "00" & x"3ba" => DATA <= x"4e73";
            when "00" & x"3bb" => DATA <= x"203c";
            when "00" & x"3bc" => DATA <= x"003f";
            when "00" & x"3bd" => DATA <= x"2dd4";
            when "00" & x"3be" => DATA <= x"207c";
            when "00" & x"3bf" => DATA <= x"0000";
            when "00" & x"3c0" => DATA <= x"002b";
            when "00" & x"3c1" => DATA <= x"4e4c";
            when "00" & x"3c2" => DATA <= x"4e75";
            when "00" & x"3c3" => DATA <= x"7000";
            when "00" & x"3c4" => DATA <= x"2a40";
            when "00" & x"3c5" => DATA <= x"206d";
            when "00" & x"3c6" => DATA <= x"000c";
            when "00" & x"3c7" => DATA <= x"43fa";
            when "00" & x"3c8" => DATA <= x"000e";
            when "00" & x"3c9" => DATA <= x"2b49";
            when "00" & x"3ca" => DATA <= x"000c";
            when "00" & x"3cb" => DATA <= x"2e0f";
            when "00" & x"3cc" => DATA <= x"2c07";
            when "00" & x"3cd" => DATA <= x"4efa";
            when "00" & x"3ce" => DATA <= x"0003";
            when "00" & x"3cf" => DATA <= x"2b48";
            when "00" & x"3d0" => DATA <= x"000c";
            when "00" & x"3d1" => DATA <= x"9e8f";
            when "00" & x"3d2" => DATA <= x"7001";
            when "00" & x"3d3" => DATA <= x"0c07";
            when "00" & x"3d4" => DATA <= x"0012";
            when "00" & x"3d5" => DATA <= x"6754";
            when "00" & x"3d6" => DATA <= x"7002";
            when "00" & x"3d7" => DATA <= x"0c07";
            when "00" & x"3d8" => DATA <= x"003e";
            when "00" & x"3d9" => DATA <= x"674c";
            when "00" & x"3da" => DATA <= x"7007";
            when "00" & x"3db" => DATA <= x"0c07";
            when "00" & x"3dc" => DATA <= x"0026";
            when "00" & x"3dd" => DATA <= x"6744";
            when "00" & x"3de" => DATA <= x"7008";
            when "00" & x"3df" => DATA <= x"0c07";
            when "00" & x"3e0" => DATA <= x"001c";
            when "00" & x"3e1" => DATA <= x"673c";
            when "00" & x"3e2" => DATA <= x"7005";
            when "00" & x"3e3" => DATA <= x"0c07";
            when "00" & x"3e4" => DATA <= x"0010";
            when "00" & x"3e5" => DATA <= x"6734";
            when "00" & x"3e6" => DATA <= x"70ff";
            when "00" & x"3e7" => DATA <= x"0c07";
            when "00" & x"3e8" => DATA <= x"0024";
            when "00" & x"3e9" => DATA <= x"662c";
            when "00" & x"3ea" => DATA <= x"206d";
            when "00" & x"3eb" => DATA <= x"001a";
            when "00" & x"3ec" => DATA <= x"226d";
            when "00" & x"3ed" => DATA <= x"007e";
            when "00" & x"3ee" => DATA <= x"45fa";
            when "00" & x"3ef" => DATA <= x"001a";
            when "00" & x"3f0" => DATA <= x"2b4a";
            when "00" & x"3f1" => DATA <= x"007e";
            when "00" & x"3f2" => DATA <= x"45fa";
            when "00" & x"3f3" => DATA <= x"0010";
            when "00" & x"3f4" => DATA <= x"2b4a";
            when "00" & x"3f5" => DATA <= x"001a";
            when "00" & x"3f6" => DATA <= x"7003";
            when "00" & x"3f7" => DATA <= x"06fa";
            when "00" & x"3f8" => DATA <= x"0000";
            when "00" & x"3f9" => DATA <= x"0002";
            when "00" & x"3fa" => DATA <= x"ffff";
            when "00" & x"3fb" => DATA <= x"7004";
            when "00" & x"3fc" => DATA <= x"2b49";
            when "00" & x"3fd" => DATA <= x"007e";
            when "00" & x"3fe" => DATA <= x"2b48";
            when "00" & x"3ff" => DATA <= x"001a";
            when "00" & x"400" => DATA <= x"2e46";
            when "00" & x"401" => DATA <= x"4e75";
            when "00" & x"402" => DATA <= x"7000";
            when "00" & x"403" => DATA <= x"2a40";
            when "00" & x"404" => DATA <= x"206d";
            when "00" & x"405" => DATA <= x"002c";
            when "00" & x"406" => DATA <= x"43fa";
            when "00" & x"407" => DATA <= x"000e";
            when "00" & x"408" => DATA <= x"2b49";
            when "00" & x"409" => DATA <= x"002c";
            when "00" & x"40a" => DATA <= x"2e0f";
            when "00" & x"40b" => DATA <= x"70ff";
            when "00" & x"40c" => DATA <= x"6000";
            when "00" & x"40d" => DATA <= x"0004";
            when "00" & x"40e" => DATA <= x"7000";
            when "00" & x"40f" => DATA <= x"2e47";
            when "00" & x"410" => DATA <= x"2b48";
            when "00" & x"411" => DATA <= x"002c";
            when "00" & x"412" => DATA <= x"4e75";
            when "00" & x"413" => DATA <= x"7000";
            when "00" & x"414" => DATA <= x"4e75";
            when "00" & x"415" => DATA <= x"13fc";
            when "00" & x"416" => DATA <= x"00f0";
            when "00" & x"417" => DATA <= x"003f";
            when "00" & x"418" => DATA <= x"0000";
            when "00" & x"419" => DATA <= x"13fc";
            when "00" & x"41a" => DATA <= x"00ff";
            when "00" & x"41b" => DATA <= x"003f";
            when "00" & x"41c" => DATA <= x"0000";
            when "00" & x"41d" => DATA <= x"4e75";
            when "00" & x"41e" => DATA <= x"13fc";
            when "00" & x"41f" => DATA <= x"00aa";
            when "00" & x"420" => DATA <= x"003f";
            when "00" & x"421" => DATA <= x"5555";
            when "00" & x"422" => DATA <= x"13fc";
            when "00" & x"423" => DATA <= x"0055";
            when "00" & x"424" => DATA <= x"003f";
            when "00" & x"425" => DATA <= x"aaaa";
            when "00" & x"426" => DATA <= x"13fc";
            when "00" & x"427" => DATA <= x"0090";
            when "00" & x"428" => DATA <= x"003f";
            when "00" & x"429" => DATA <= x"5555";
            when "00" & x"42a" => DATA <= x"13c0";
            when "00" & x"42b" => DATA <= x"003f";
            when "00" & x"42c" => DATA <= x"0000";
            when "00" & x"42d" => DATA <= x"e140";
            when "00" & x"42e" => DATA <= x"61cc";
            when "00" & x"42f" => DATA <= x"13fc";
            when "00" & x"430" => DATA <= x"00aa";
            when "00" & x"431" => DATA <= x"003f";
            when "00" & x"432" => DATA <= x"5555";
            when "00" & x"433" => DATA <= x"13fc";
            when "00" & x"434" => DATA <= x"0055";
            when "00" & x"435" => DATA <= x"003f";
            when "00" & x"436" => DATA <= x"aaaa";
            when "00" & x"437" => DATA <= x"13fc";
            when "00" & x"438" => DATA <= x"0090";
            when "00" & x"439" => DATA <= x"003f";
            when "00" & x"43a" => DATA <= x"5555";
            when "00" & x"43b" => DATA <= x"13c0";
            when "00" & x"43c" => DATA <= x"003f";
            when "00" & x"43d" => DATA <= x"0001";
            when "00" & x"43e" => DATA <= x"61ac";
            when "00" & x"43f" => DATA <= x"4e75";
            when "00" & x"440" => DATA <= x"be3c";
            when "00" & x"441" => DATA <= x"0008";
            when "00" & x"442" => DATA <= x"6400";
            when "00" & x"443" => DATA <= x"0012";
            when "00" & x"444" => DATA <= x"e147";
            when "00" & x"445" => DATA <= x"e147";
            when "00" & x"446" => DATA <= x"223c";
            when "00" & x"447" => DATA <= x"0000";
            when "00" & x"448" => DATA <= x"ffff";
            when "00" & x"449" => DATA <= x"1015";
            when "00" & x"44a" => DATA <= x"6100";
            when "00" & x"44b" => DATA <= x"0004";
            when "00" & x"44c" => DATA <= x"4e75";
            when "00" & x"44d" => DATA <= x"b016";
            when "00" & x"44e" => DATA <= x"6700";
            when "00" & x"44f" => DATA <= x"0026";
            when "00" & x"450" => DATA <= x"13fc";
            when "00" & x"451" => DATA <= x"00aa";
            when "00" & x"452" => DATA <= x"003f";
            when "00" & x"453" => DATA <= x"5555";
            when "00" & x"454" => DATA <= x"13fc";
            when "00" & x"455" => DATA <= x"0055";
            when "00" & x"456" => DATA <= x"003f";
            when "00" & x"457" => DATA <= x"aaaa";
            when "00" & x"458" => DATA <= x"13fc";
            when "00" & x"459" => DATA <= x"00a0";
            when "00" & x"45a" => DATA <= x"003f";
            when "00" & x"45b" => DATA <= x"5555";
            when "00" & x"45c" => DATA <= x"1016";
            when "00" & x"45d" => DATA <= x"0c16";
            when "00" & x"45e" => DATA <= x"0002";
            when "00" & x"45f" => DATA <= x"66fa";
            when "00" & x"460" => DATA <= x"6100";
            when "00" & x"461" => DATA <= x"ff68";
            when "00" & x"462" => DATA <= x"4e75";
            when "00" & x"463" => DATA <= x"2f08";
            when "00" & x"464" => DATA <= x"2f38";
            when "00" & x"465" => DATA <= x"0000";
            when "00" & x"466" => DATA <= x"207c";
            when "00" & x"467" => DATA <= x"0000";
            when "00" & x"468" => DATA <= x"0000";
            when "00" & x"469" => DATA <= x"21fc";
            when "00" & x"46a" => DATA <= x"dead";
            when "00" & x"46b" => DATA <= x"beef";
            when "00" & x"46c" => DATA <= x"0000";
            when "00" & x"46d" => DATA <= x"d1fc";
            when "00" & x"46e" => DATA <= x"0000";
            when "00" & x"46f" => DATA <= x"0400";
            when "00" & x"470" => DATA <= x"0c90";
            when "00" & x"471" => DATA <= x"dead";
            when "00" & x"472" => DATA <= x"beef";
            when "00" & x"473" => DATA <= x"6700";
            when "00" & x"474" => DATA <= x"000a";
            when "00" & x"475" => DATA <= x"b1fc";
            when "00" & x"476" => DATA <= x"0030";
            when "00" & x"477" => DATA <= x"0000";
            when "00" & x"478" => DATA <= x"65e8";
            when "00" & x"479" => DATA <= x"2008";
            when "00" & x"47a" => DATA <= x"21df";
            when "00" & x"47b" => DATA <= x"0000";
            when "00" & x"47c" => DATA <= x"205f";
            when "00" & x"47d" => DATA <= x"4e75";
            when "00" & x"47e" => DATA <= x"2f0e";
            when "00" & x"47f" => DATA <= x"2f09";
            when "00" & x"480" => DATA <= x"2f08";
            when "00" & x"481" => DATA <= x"2f01";
            when "00" & x"482" => DATA <= x"c188";
            when "00" & x"483" => DATA <= x"0280";
            when "00" & x"484" => DATA <= x"00fd";
            when "00" & x"485" => DATA <= x"ffff";
            when "00" & x"486" => DATA <= x"43f9";
            when "00" & x"487" => DATA <= x"003f";
            when "00" & x"488" => DATA <= x"2f50";
            when "00" & x"489" => DATA <= x"b099";
            when "00" & x"48a" => DATA <= x"6700";
            when "00" & x"48b" => DATA <= x"0014";
            when "00" & x"48c" => DATA <= x"2219";
            when "00" & x"48d" => DATA <= x"b23c";
            when "00" & x"48e" => DATA <= x"00ff";
            when "00" & x"48f" => DATA <= x"6700";
            when "00" & x"490" => DATA <= x"0082";
            when "00" & x"491" => DATA <= x"b23c";
            when "00" & x"492" => DATA <= x"0000";
            when "00" & x"493" => DATA <= x"66f0";
            when "00" & x"494" => DATA <= x"60e8";
            when "00" & x"495" => DATA <= x"2c59";
            when "00" & x"496" => DATA <= x"c188";
            when "00" & x"497" => DATA <= x"bdfc";
            when "00" & x"498" => DATA <= x"0000";
            when "00" & x"499" => DATA <= x"0504";
            when "00" & x"49a" => DATA <= x"6400";
            when "00" & x"49b" => DATA <= x"0004";
            when "00" & x"49c" => DATA <= x"2c56";
            when "00" & x"49d" => DATA <= x"221f";
            when "00" & x"49e" => DATA <= x"205f";
            when "00" & x"49f" => DATA <= x"225f";
            when "00" & x"4a0" => DATA <= x"4e96";
            when "00" & x"4a1" => DATA <= x"6900";
            when "00" & x"4a2" => DATA <= x"001a";
            when "00" & x"4a3" => DATA <= x"6500";
            when "00" & x"4a4" => DATA <= x"000a";
            when "00" & x"4a5" => DATA <= x"2c5f";
            when "00" & x"4a6" => DATA <= x"0257";
            when "00" & x"4a7" => DATA <= x"fffc";
            when "00" & x"4a8" => DATA <= x"4e73";
            when "00" & x"4a9" => DATA <= x"2c5f";
            when "00" & x"4aa" => DATA <= x"0257";
            when "00" & x"4ab" => DATA <= x"fffd";
            when "00" & x"4ac" => DATA <= x"0057";
            when "00" & x"4ad" => DATA <= x"0001";
            when "00" & x"4ae" => DATA <= x"4e73";
            when "00" & x"4af" => DATA <= x"6500";
            when "00" & x"4b0" => DATA <= x"000e";
            when "00" & x"4b1" => DATA <= x"0057";
            when "00" & x"4b2" => DATA <= x"0002";
            when "00" & x"4b3" => DATA <= x"0257";
            when "00" & x"4b4" => DATA <= x"fffe";
            when "00" & x"4b5" => DATA <= x"6000";
            when "00" & x"4b6" => DATA <= x"0006";
            when "00" & x"4b7" => DATA <= x"0057";
            when "00" & x"4b8" => DATA <= x"0003";
            when "00" & x"4b9" => DATA <= x"2c5f";
            when "00" & x"4ba" => DATA <= x"c188";
            when "00" & x"4bb" => DATA <= x"0800";
            when "00" & x"4bc" => DATA <= x"0011";
            when "00" & x"4bd" => DATA <= x"6700";
            when "00" & x"4be" => DATA <= x"0006";
            when "00" & x"4bf" => DATA <= x"c188";
            when "00" & x"4c0" => DATA <= x"4e73";
            when "00" & x"4c1" => DATA <= x"c188";
            when "00" & x"4c2" => DATA <= x"2f01";
            when "00" & x"4c3" => DATA <= x"7206";
            when "00" & x"4c4" => DATA <= x"6100";
            when "00" & x"4c5" => DATA <= x"07c6";
            when "00" & x"4c6" => DATA <= x"221f";
            when "00" & x"4c7" => DATA <= x"21c0";
            when "00" & x"4c8" => DATA <= x"0514";
            when "00" & x"4c9" => DATA <= x"21ef";
            when "00" & x"4ca" => DATA <= x"0002";
            when "00" & x"4cb" => DATA <= x"0510";
            when "00" & x"4cc" => DATA <= x"2f79";
            when "00" & x"4cd" => DATA <= x"0000";
            when "00" & x"4ce" => DATA <= x"0404";
            when "00" & x"4cf" => DATA <= x"0002";
            when "00" & x"4d0" => DATA <= x"4e73";
            when "00" & x"4d1" => DATA <= x"221f";
            when "00" & x"4d2" => DATA <= x"205f";
            when "00" & x"4d3" => DATA <= x"225f";
            when "00" & x"4d4" => DATA <= x"2040";
            when "00" & x"4d5" => DATA <= x"c0bc";
            when "00" & x"4d6" => DATA <= x"00fd";
            when "00" & x"4d7" => DATA <= x"ff00";
            when "00" & x"4d8" => DATA <= x"b0bc";
            when "00" & x"4d9" => DATA <= x"0000";
            when "00" & x"4da" => DATA <= x"0100";
            when "00" & x"4db" => DATA <= x"6600";
            when "00" & x"4dc" => DATA <= x"0012";
            when "00" & x"4dd" => DATA <= x"2008";
            when "00" & x"4de" => DATA <= x"4eb9";
            when "00" & x"4df" => DATA <= x"003f";
            when "00" & x"4e0" => DATA <= x"09e0";
            when "00" & x"4e1" => DATA <= x"2c5f";
            when "00" & x"4e2" => DATA <= x"0257";
            when "00" & x"4e3" => DATA <= x"fffc";
            when "00" & x"4e4" => DATA <= x"4e73";
            when "00" & x"4e5" => DATA <= x"2008";
            when "00" & x"4e6" => DATA <= x"2c78";
            when "00" & x"4e7" => DATA <= x"0460";
            when "00" & x"4e8" => DATA <= x"21ef";
            when "00" & x"4e9" => DATA <= x"0006";
            when "00" & x"4ea" => DATA <= x"0510";
            when "00" & x"4eb" => DATA <= x"4e96";
            when "00" & x"4ec" => DATA <= x"2c5f";
            when "00" & x"4ed" => DATA <= x"0057";
            when "00" & x"4ee" => DATA <= x"0002";
            when "00" & x"4ef" => DATA <= x"4e73";
            when "00" & x"4f0" => DATA <= x"201f";
            when "00" & x"4f1" => DATA <= x"6000";
            when "00" & x"4f2" => DATA <= x"0002";
            when "00" & x"4f3" => DATA <= x"2f38";
            when "00" & x"4f4" => DATA <= x"040c";
            when "00" & x"4f5" => DATA <= x"4e75";
            when "00" & x"4f6" => DATA <= x"2f00";
            when "00" & x"4f7" => DATA <= x"202f";
            when "00" & x"4f8" => DATA <= x"0004";
            when "00" & x"4f9" => DATA <= x"6100";
            when "00" & x"4fa" => DATA <= x"000a";
            when "00" & x"4fb" => DATA <= x"2f40";
            when "00" & x"4fc" => DATA <= x"0004";
            when "00" & x"4fd" => DATA <= x"201f";
            when "00" & x"4fe" => DATA <= x"4e75";
            when "00" & x"4ff" => DATA <= x"2f08";
            when "00" & x"500" => DATA <= x"2040";
            when "00" & x"501" => DATA <= x"1018";
            when "00" & x"502" => DATA <= x"6700";
            when "00" & x"503" => DATA <= x"0006";
            when "00" & x"504" => DATA <= x"61dc";
            when "00" & x"505" => DATA <= x"60f6";
            when "00" & x"506" => DATA <= x"2008";
            when "00" & x"507" => DATA <= x"205f";
            when "00" & x"508" => DATA <= x"4e75";
            when "00" & x"509" => DATA <= x"2f00";
            when "00" & x"50a" => DATA <= x"700a";
            when "00" & x"50b" => DATA <= x"61ce";
            when "00" & x"50c" => DATA <= x"700d";
            when "00" & x"50d" => DATA <= x"61ca";
            when "00" & x"50e" => DATA <= x"201f";
            when "00" & x"50f" => DATA <= x"4e75";
            when "00" & x"510" => DATA <= x"7000";
            when "00" & x"511" => DATA <= x"6100";
            when "00" & x"512" => DATA <= x"f9be";
            when "00" & x"513" => DATA <= x"6100";
            when "00" & x"514" => DATA <= x"f9a8";
            when "00" & x"515" => DATA <= x"e000";
            when "00" & x"516" => DATA <= x"6000";
            when "00" & x"517" => DATA <= x"f9a2";
            when "00" & x"518" => DATA <= x"2f0e";
            when "00" & x"519" => DATA <= x"2f00";
            when "00" & x"51a" => DATA <= x"2c40";
            when "00" & x"51b" => DATA <= x"6100";
            when "00" & x"51c" => DATA <= x"1ce8";
            when "00" & x"51d" => DATA <= x"101e";
            when "00" & x"51e" => DATA <= x"b03c";
            when "00" & x"51f" => DATA <= x"002a";
            when "00" & x"520" => DATA <= x"67f4";
            when "00" & x"521" => DATA <= x"1026";
            when "00" & x"522" => DATA <= x"43f9";
            when "00" & x"523" => DATA <= x"003f";
            when "00" & x"524" => DATA <= x"35cc";
            when "00" & x"525" => DATA <= x"2f0e";
            when "00" & x"526" => DATA <= x"2459";
            when "00" & x"527" => DATA <= x"b4fc";
            when "00" & x"528" => DATA <= x"ffff";
            when "00" & x"529" => DATA <= x"6700";
            when "00" & x"52a" => DATA <= x"0050";
            when "00" & x"52b" => DATA <= x"101e";
            when "00" & x"52c" => DATA <= x"0200";
            when "00" & x"52d" => DATA <= x"00df";
            when "00" & x"52e" => DATA <= x"b019";
            when "00" & x"52f" => DATA <= x"6600";
            when "00" & x"530" => DATA <= x"003a";
            when "00" & x"531" => DATA <= x"0c16";
            when "00" & x"532" => DATA <= x"002e";
            when "00" & x"533" => DATA <= x"6700";
            when "00" & x"534" => DATA <= x"0010";
            when "00" & x"535" => DATA <= x"0c11";
            when "00" & x"536" => DATA <= x"0020";
            when "00" & x"537" => DATA <= x"6700";
            when "00" & x"538" => DATA <= x"0008";
            when "00" & x"539" => DATA <= x"0c11";
            when "00" & x"53a" => DATA <= x"0000";
            when "00" & x"53b" => DATA <= x"66de";
            when "00" & x"53c" => DATA <= x"0c16";
            when "00" & x"53d" => DATA <= x"000d";
            when "00" & x"53e" => DATA <= x"6700";
            when "00" & x"53f" => DATA <= x"000a";
            when "00" & x"540" => DATA <= x"0c16";
            when "00" & x"541" => DATA <= x"0020";
            when "00" & x"542" => DATA <= x"6600";
            when "00" & x"543" => DATA <= x"0014";
            when "00" & x"544" => DATA <= x"6100";
            when "00" & x"545" => DATA <= x"1c96";
            when "00" & x"546" => DATA <= x"225f";
            when "00" & x"547" => DATA <= x"4e92";
            when "00" & x"548" => DATA <= x"201f";
            when "00" & x"549" => DATA <= x"2c5f";
            when "00" & x"54a" => DATA <= x"6500";
            when "00" & x"54b" => DATA <= x"0012";
            when "00" & x"54c" => DATA <= x"4e75";
            when "00" & x"54d" => DATA <= x"0c19";
            when "00" & x"54e" => DATA <= x"0000";
            when "00" & x"54f" => DATA <= x"66fa";
            when "00" & x"550" => DATA <= x"2c5f";
            when "00" & x"551" => DATA <= x"60a6";
            when "00" & x"552" => DATA <= x"2c5f";
            when "00" & x"553" => DATA <= x"201f";
            when "00" & x"554" => DATA <= x"2f01";
            when "00" & x"555" => DATA <= x"7204";
            when "00" & x"556" => DATA <= x"6100";
            when "00" & x"557" => DATA <= x"06a2";
            when "00" & x"558" => DATA <= x"221f";
            when "00" & x"559" => DATA <= x"2c40";
            when "00" & x"55a" => DATA <= x"7002";
            when "00" & x"55b" => DATA <= x"6100";
            when "00" & x"55c" => DATA <= x"f92a";
            when "00" & x"55d" => DATA <= x"6100";
            when "00" & x"55e" => DATA <= x"f97a";
            when "00" & x"55f" => DATA <= x"6100";
            when "00" & x"560" => DATA <= x"f910";
            when "00" & x"561" => DATA <= x"2c5f";
            when "00" & x"562" => DATA <= x"b03c";
            when "00" & x"563" => DATA <= x"0080";
            when "00" & x"564" => DATA <= x"6700";
            when "00" & x"565" => DATA <= x"00b6";
            when "00" & x"566" => DATA <= x"023c";
            when "00" & x"567" => DATA <= x"00fd";
            when "00" & x"568" => DATA <= x"4e75";
            when "00" & x"569" => DATA <= x"b03c";
            when "00" & x"56a" => DATA <= x"0080";
            when "00" & x"56b" => DATA <= x"6400";
            when "00" & x"56c" => DATA <= x"002a";
            when "00" & x"56d" => DATA <= x"b03c";
            when "00" & x"56e" => DATA <= x"007e";
            when "00" & x"56f" => DATA <= x"6600";
            when "00" & x"570" => DATA <= x"0002";
            when "00" & x"571" => DATA <= x"2f00";
            when "00" & x"572" => DATA <= x"103c";
            when "00" & x"573" => DATA <= x"0004";
            when "00" & x"574" => DATA <= x"6100";
            when "00" & x"575" => DATA <= x"f8f8";
            when "00" & x"576" => DATA <= x"1001";
            when "00" & x"577" => DATA <= x"6100";
            when "00" & x"578" => DATA <= x"f8f2";
            when "00" & x"579" => DATA <= x"2017";
            when "00" & x"57a" => DATA <= x"6100";
            when "00" & x"57b" => DATA <= x"f8ec";
            when "00" & x"57c" => DATA <= x"6100";
            when "00" & x"57d" => DATA <= x"f8d6";
            when "00" & x"57e" => DATA <= x"1200";
            when "00" & x"57f" => DATA <= x"201f";
            when "00" & x"580" => DATA <= x"4e75";
            when "00" & x"581" => DATA <= x"b03c";
            when "00" & x"582" => DATA <= x"0082";
            when "00" & x"583" => DATA <= x"6700";
            when "00" & x"584" => DATA <= x"005a";
            when "00" & x"585" => DATA <= x"b03c";
            when "00" & x"586" => DATA <= x"0083";
            when "00" & x"587" => DATA <= x"6700";
            when "00" & x"588" => DATA <= x"005c";
            when "00" & x"589" => DATA <= x"b03c";
            when "00" & x"58a" => DATA <= x"0084";
            when "00" & x"58b" => DATA <= x"6700";
            when "00" & x"58c" => DATA <= x"005e";
            when "00" & x"58d" => DATA <= x"2f00";
            when "00" & x"58e" => DATA <= x"103c";
            when "00" & x"58f" => DATA <= x"0006";
            when "00" & x"590" => DATA <= x"6100";
            when "00" & x"591" => DATA <= x"f8c0";
            when "00" & x"592" => DATA <= x"1001";
            when "00" & x"593" => DATA <= x"6100";
            when "00" & x"594" => DATA <= x"f8ba";
            when "00" & x"595" => DATA <= x"1002";
            when "00" & x"596" => DATA <= x"6100";
            when "00" & x"597" => DATA <= x"f8b4";
            when "00" & x"598" => DATA <= x"201f";
            when "00" & x"599" => DATA <= x"6100";
            when "00" & x"59a" => DATA <= x"f8ae";
            when "00" & x"59b" => DATA <= x"b03c";
            when "00" & x"59c" => DATA <= x"008e";
            when "00" & x"59d" => DATA <= x"6700";
            when "00" & x"59e" => DATA <= x"0044";
            when "00" & x"59f" => DATA <= x"b03c";
            when "00" & x"5a0" => DATA <= x"009d";
            when "00" & x"5a1" => DATA <= x"6700";
            when "00" & x"5a2" => DATA <= x"009e";
            when "00" & x"5a3" => DATA <= x"2f00";
            when "00" & x"5a4" => DATA <= x"6100";
            when "00" & x"5a5" => DATA <= x"f886";
            when "00" & x"5a6" => DATA <= x"3f00";
            when "00" & x"5a7" => DATA <= x"6100";
            when "00" & x"5a8" => DATA <= x"f880";
            when "00" & x"5a9" => DATA <= x"1400";
            when "00" & x"5aa" => DATA <= x"6100";
            when "00" & x"5ab" => DATA <= x"f87a";
            when "00" & x"5ac" => DATA <= x"1200";
            when "00" & x"5ad" => DATA <= x"201f";
            when "00" & x"5ae" => DATA <= x"e000";
            when "00" & x"5af" => DATA <= x"201f";
            when "00" & x"5b0" => DATA <= x"4e75";
            when "00" & x"5b1" => DATA <= x"3238";
            when "00" & x"5b2" => DATA <= x"0524";
            when "00" & x"5b3" => DATA <= x"2401";
            when "00" & x"5b4" => DATA <= x"e082";
            when "00" & x"5b5" => DATA <= x"4e75";
            when "00" & x"5b6" => DATA <= x"2238";
            when "00" & x"5b7" => DATA <= x"0504";
            when "00" & x"5b8" => DATA <= x"2401";
            when "00" & x"5b9" => DATA <= x"e082";
            when "00" & x"5ba" => DATA <= x"4e75";
            when "00" & x"5bb" => DATA <= x"2238";
            when "00" & x"5bc" => DATA <= x"0500";
            when "00" & x"5bd" => DATA <= x"2401";
            when "00" & x"5be" => DATA <= x"e082";
            when "00" & x"5bf" => DATA <= x"4e75";
            when "00" & x"5c0" => DATA <= x"2c78";
            when "00" & x"5c1" => DATA <= x"0520";
            when "00" & x"5c2" => DATA <= x"122e";
            when "00" & x"5c3" => DATA <= x"0006";
            when "00" & x"5c4" => DATA <= x"7000";
            when "00" & x"5c5" => DATA <= x"102e";
            when "00" & x"5c6" => DATA <= x"0007";
            when "00" & x"5c7" => DATA <= x"ddc0";
            when "00" & x"5c8" => DATA <= x"4a1e";
            when "00" & x"5c9" => DATA <= x"6600";
            when "00" & x"5ca" => DATA <= x"0026";
            when "00" & x"5cb" => DATA <= x"0c1e";
            when "00" & x"5cc" => DATA <= x"0028";
            when "00" & x"5cd" => DATA <= x"6600";
            when "00" & x"5ce" => DATA <= x"001e";
            when "00" & x"5cf" => DATA <= x"0c1e";
            when "00" & x"5d0" => DATA <= x"0043";
            when "00" & x"5d1" => DATA <= x"6600";
            when "00" & x"5d2" => DATA <= x"0016";
            when "00" & x"5d3" => DATA <= x"0c1e";
            when "00" & x"5d4" => DATA <= x"0029";
            when "00" & x"5d5" => DATA <= x"6600";
            when "00" & x"5d6" => DATA <= x"000e";
            when "00" & x"5d7" => DATA <= x"0201";
            when "00" & x"5d8" => DATA <= x"000f";
            when "00" & x"5d9" => DATA <= x"0c01";
            when "00" & x"5da" => DATA <= x"0003";
            when "00" & x"5db" => DATA <= x"6600";
            when "00" & x"5dc" => DATA <= x"0018";
            when "00" & x"5dd" => DATA <= x"2c78";
            when "00" & x"5de" => DATA <= x"0520";
            when "00" & x"5df" => DATA <= x"7001";
            when "00" & x"5e0" => DATA <= x"223c";
            when "00" & x"5e1" => DATA <= x"0000";
            when "00" & x"5e2" => DATA <= x"052d";
            when "00" & x"5e3" => DATA <= x"6100";
            when "00" & x"5e4" => DATA <= x"001c";
            when "00" & x"5e5" => DATA <= x"7001";
            when "00" & x"5e6" => DATA <= x"4ed6";
            when "00" & x"5e7" => DATA <= x"4e75";
            when "00" & x"5e8" => DATA <= x"203c";
            when "00" & x"5e9" => DATA <= x"003f";
            when "00" & x"5ea" => DATA <= x"2da0";
            when "00" & x"5eb" => DATA <= x"21fc";
            when "00" & x"5ec" => DATA <= x"0000";
            when "00" & x"5ed" => DATA <= x"0000";
            when "00" & x"5ee" => DATA <= x"0510";
            when "00" & x"5ef" => DATA <= x"6000";
            when "00" & x"5f0" => DATA <= x"0540";
            when "00" & x"5f1" => DATA <= x"4e75";
            when "00" & x"5f2" => DATA <= x"b0bc";
            when "00" & x"5f3" => DATA <= x"0000";
            when "00" & x"5f4" => DATA <= x"00ff";
            when "00" & x"5f5" => DATA <= x"6200";
            when "00" & x"5f6" => DATA <= x"00d8";
            when "00" & x"5f7" => DATA <= x"2f0e";
            when "00" & x"5f8" => DATA <= x"2f00";
            when "00" & x"5f9" => DATA <= x"2f01";
            when "00" & x"5fa" => DATA <= x"2f02";
            when "00" & x"5fb" => DATA <= x"2c41";
            when "00" & x"5fc" => DATA <= x"4a40";
            when "00" & x"5fd" => DATA <= x"6600";
            when "00" & x"5fe" => DATA <= x"003c";
            when "00" & x"5ff" => DATA <= x"2f03";
            when "00" & x"600" => DATA <= x"2f04";
            when "00" & x"601" => DATA <= x"3038";
            when "00" & x"602" => DATA <= x"0524";
            when "00" & x"603" => DATA <= x"4840";
            when "00" & x"604" => DATA <= x"3016";
            when "00" & x"605" => DATA <= x"7200";
            when "00" & x"606" => DATA <= x"122e";
            when "00" & x"607" => DATA <= x"0002";
            when "00" & x"608" => DATA <= x"7400";
            when "00" & x"609" => DATA <= x"142e";
            when "00" & x"60a" => DATA <= x"0003";
            when "00" & x"60b" => DATA <= x"7600";
            when "00" & x"60c" => DATA <= x"162e";
            when "00" & x"60d" => DATA <= x"0004";
            when "00" & x"60e" => DATA <= x"7800";
            when "00" & x"60f" => DATA <= x"6100";
            when "00" & x"610" => DATA <= x"08cc";
            when "00" & x"611" => DATA <= x"281f";
            when "00" & x"612" => DATA <= x"261f";
            when "00" & x"613" => DATA <= x"241f";
            when "00" & x"614" => DATA <= x"2401";
            when "00" & x"615" => DATA <= x"5242";
            when "00" & x"616" => DATA <= x"221f";
            when "00" & x"617" => DATA <= x"201f";
            when "00" & x"618" => DATA <= x"2c5f";
            when "00" & x"619" => DATA <= x"023c";
            when "00" & x"61a" => DATA <= x"00fd";
            when "00" & x"61b" => DATA <= x"4e75";
            when "00" & x"61c" => DATA <= x"7200";
            when "00" & x"61d" => DATA <= x"7400";
            when "00" & x"61e" => DATA <= x"b03c";
            when "00" & x"61f" => DATA <= x"0014";
            when "00" & x"620" => DATA <= x"6200";
            when "00" & x"621" => DATA <= x"001e";
            when "00" & x"622" => DATA <= x"207c";
            when "00" & x"623" => DATA <= x"003f";
            when "00" & x"624" => DATA <= x"2f28";
            when "00" & x"625" => DATA <= x"d1c0";
            when "00" & x"626" => DATA <= x"5348";
            when "00" & x"627" => DATA <= x"1210";
            when "00" & x"628" => DATA <= x"207c";
            when "00" & x"629" => DATA <= x"003f";
            when "00" & x"62a" => DATA <= x"2f3c";
            when "00" & x"62b" => DATA <= x"d1c0";
            when "00" & x"62c" => DATA <= x"5348";
            when "00" & x"62d" => DATA <= x"1410";
            when "00" & x"62e" => DATA <= x"6000";
            when "00" & x"62f" => DATA <= x"0018";
            when "00" & x"630" => DATA <= x"b03c";
            when "00" & x"631" => DATA <= x"007f";
            when "00" & x"632" => DATA <= x"6200";
            when "00" & x"633" => DATA <= x"000a";
            when "00" & x"634" => DATA <= x"7210";
            when "00" & x"635" => DATA <= x"7410";
            when "00" & x"636" => DATA <= x"6000";
            when "00" & x"637" => DATA <= x"0008";
            when "00" & x"638" => DATA <= x"1216";
            when "00" & x"639" => DATA <= x"142e";
            when "00" & x"63a" => DATA <= x"0001";
            when "00" & x"63b" => DATA <= x"2f00";
            when "00" & x"63c" => DATA <= x"103c";
            when "00" & x"63d" => DATA <= x"0008";
            when "00" & x"63e" => DATA <= x"6100";
            when "00" & x"63f" => DATA <= x"f764";
            when "00" & x"640" => DATA <= x"201f";
            when "00" & x"641" => DATA <= x"6100";
            when "00" & x"642" => DATA <= x"f75e";
            when "00" & x"643" => DATA <= x"1001";
            when "00" & x"644" => DATA <= x"6100";
            when "00" & x"645" => DATA <= x"f758";
            when "00" & x"646" => DATA <= x"5341";
            when "00" & x"647" => DATA <= x"6b00";
            when "00" & x"648" => DATA <= x"000e";
            when "00" & x"649" => DATA <= x"1036";
            when "00" & x"64a" => DATA <= x"1000";
            when "00" & x"64b" => DATA <= x"6100";
            when "00" & x"64c" => DATA <= x"f74a";
            when "00" & x"64d" => DATA <= x"51c9";
            when "00" & x"64e" => DATA <= x"fff6";
            when "00" & x"64f" => DATA <= x"1002";
            when "00" & x"650" => DATA <= x"6100";
            when "00" & x"651" => DATA <= x"f740";
            when "00" & x"652" => DATA <= x"5342";
            when "00" & x"653" => DATA <= x"6b00";
            when "00" & x"654" => DATA <= x"000e";
            when "00" & x"655" => DATA <= x"6100";
            when "00" & x"656" => DATA <= x"f724";
            when "00" & x"657" => DATA <= x"1d80";
            when "00" & x"658" => DATA <= x"2000";
            when "00" & x"659" => DATA <= x"51ca";
            when "00" & x"65a" => DATA <= x"fff6";
            when "00" & x"65b" => DATA <= x"241f";
            when "00" & x"65c" => DATA <= x"221f";
            when "00" & x"65d" => DATA <= x"201f";
            when "00" & x"65e" => DATA <= x"2c5f";
            when "00" & x"65f" => DATA <= x"023c";
            when "00" & x"660" => DATA <= x"00fd";
            when "00" & x"661" => DATA <= x"4e75";
            when "00" & x"662" => DATA <= x"003c";
            when "00" & x"663" => DATA <= x"0002";
            when "00" & x"664" => DATA <= x"4e75";
            when "00" & x"665" => DATA <= x"2f00";
            when "00" & x"666" => DATA <= x"103c";
            when "00" & x"667" => DATA <= x"0014";
            when "00" & x"668" => DATA <= x"6100";
            when "00" & x"669" => DATA <= x"f710";
            when "00" & x"66a" => DATA <= x"2005";
            when "00" & x"66b" => DATA <= x"6100";
            when "00" & x"66c" => DATA <= x"f73e";
            when "00" & x"66d" => DATA <= x"2004";
            when "00" & x"66e" => DATA <= x"6100";
            when "00" & x"66f" => DATA <= x"f738";
            when "00" & x"670" => DATA <= x"2003";
            when "00" & x"671" => DATA <= x"6100";
            when "00" & x"672" => DATA <= x"f732";
            when "00" & x"673" => DATA <= x"2002";
            when "00" & x"674" => DATA <= x"6100";
            when "00" & x"675" => DATA <= x"f72c";
            when "00" & x"676" => DATA <= x"2c41";
            when "00" & x"677" => DATA <= x"6100";
            when "00" & x"678" => DATA <= x"f746";
            when "00" & x"679" => DATA <= x"201f";
            when "00" & x"67a" => DATA <= x"6100";
            when "00" & x"67b" => DATA <= x"f6ec";
            when "00" & x"67c" => DATA <= x"6100";
            when "00" & x"67d" => DATA <= x"f6d6";
            when "00" & x"67e" => DATA <= x"2f00";
            when "00" & x"67f" => DATA <= x"6100";
            when "00" & x"680" => DATA <= x"f706";
            when "00" & x"681" => DATA <= x"2a00";
            when "00" & x"682" => DATA <= x"6100";
            when "00" & x"683" => DATA <= x"f700";
            when "00" & x"684" => DATA <= x"2800";
            when "00" & x"685" => DATA <= x"6100";
            when "00" & x"686" => DATA <= x"f6fa";
            when "00" & x"687" => DATA <= x"2600";
            when "00" & x"688" => DATA <= x"6100";
            when "00" & x"689" => DATA <= x"f6f4";
            when "00" & x"68a" => DATA <= x"2400";
            when "00" & x"68b" => DATA <= x"201f";
            when "00" & x"68c" => DATA <= x"4e75";
            when "00" & x"68d" => DATA <= x"2f00";
            when "00" & x"68e" => DATA <= x"103c";
            when "00" & x"68f" => DATA <= x"000c";
            when "00" & x"690" => DATA <= x"6100";
            when "00" & x"691" => DATA <= x"f6c0";
            when "00" & x"692" => DATA <= x"1001";
            when "00" & x"693" => DATA <= x"6100";
            when "00" & x"694" => DATA <= x"f6ba";
            when "00" & x"695" => DATA <= x"2002";
            when "00" & x"696" => DATA <= x"6100";
            when "00" & x"697" => DATA <= x"f6e8";
            when "00" & x"698" => DATA <= x"201f";
            when "00" & x"699" => DATA <= x"6100";
            when "00" & x"69a" => DATA <= x"f6ae";
            when "00" & x"69b" => DATA <= x"6100";
            when "00" & x"69c" => DATA <= x"f698";
            when "00" & x"69d" => DATA <= x"2f00";
            when "00" & x"69e" => DATA <= x"6100";
            when "00" & x"69f" => DATA <= x"f6c8";
            when "00" & x"6a0" => DATA <= x"2400";
            when "00" & x"6a1" => DATA <= x"201f";
            when "00" & x"6a2" => DATA <= x"4e75";
            when "00" & x"6a3" => DATA <= x"103c";
            when "00" & x"6a4" => DATA <= x"000e";
            when "00" & x"6a5" => DATA <= x"4eb9";
            when "00" & x"6a6" => DATA <= x"003f";
            when "00" & x"6a7" => DATA <= x"03e2";
            when "00" & x"6a8" => DATA <= x"1001";
            when "00" & x"6a9" => DATA <= x"4eb9";
            when "00" & x"6aa" => DATA <= x"003f";
            when "00" & x"6ab" => DATA <= x"03e2";
            when "00" & x"6ac" => DATA <= x"6000";
            when "00" & x"6ad" => DATA <= x"fccc";
            when "00" & x"6ae" => DATA <= x"2f00";
            when "00" & x"6af" => DATA <= x"103c";
            when "00" & x"6b0" => DATA <= x"0010";
            when "00" & x"6b1" => DATA <= x"6100";
            when "00" & x"6b2" => DATA <= x"f67e";
            when "00" & x"6b3" => DATA <= x"1001";
            when "00" & x"6b4" => DATA <= x"6100";
            when "00" & x"6b5" => DATA <= x"f678";
            when "00" & x"6b6" => DATA <= x"2017";
            when "00" & x"6b7" => DATA <= x"6100";
            when "00" & x"6b8" => DATA <= x"f672";
            when "00" & x"6b9" => DATA <= x"6100";
            when "00" & x"6ba" => DATA <= x"f65c";
            when "00" & x"6bb" => DATA <= x"201f";
            when "00" & x"6bc" => DATA <= x"4e75";
            when "00" & x"6bd" => DATA <= x"2f00";
            when "00" & x"6be" => DATA <= x"103c";
            when "00" & x"6bf" => DATA <= x"0016";
            when "00" & x"6c0" => DATA <= x"6100";
            when "00" & x"6c1" => DATA <= x"f660";
            when "00" & x"6c2" => DATA <= x"2004";
            when "00" & x"6c3" => DATA <= x"6100";
            when "00" & x"6c4" => DATA <= x"f68e";
            when "00" & x"6c5" => DATA <= x"2003";
            when "00" & x"6c6" => DATA <= x"6100";
            when "00" & x"6c7" => DATA <= x"f688";
            when "00" & x"6c8" => DATA <= x"2002";
            when "00" & x"6c9" => DATA <= x"6100";
            when "00" & x"6ca" => DATA <= x"f682";
            when "00" & x"6cb" => DATA <= x"2001";
            when "00" & x"6cc" => DATA <= x"6100";
            when "00" & x"6cd" => DATA <= x"f648";
            when "00" & x"6ce" => DATA <= x"201f";
            when "00" & x"6cf" => DATA <= x"6100";
            when "00" & x"6d0" => DATA <= x"f676";
            when "00" & x"6d1" => DATA <= x"6100";
            when "00" & x"6d2" => DATA <= x"f62c";
            when "00" & x"6d3" => DATA <= x"2800";
            when "00" & x"6d4" => DATA <= x"6100";
            when "00" & x"6d5" => DATA <= x"f65c";
            when "00" & x"6d6" => DATA <= x"2600";
            when "00" & x"6d7" => DATA <= x"6100";
            when "00" & x"6d8" => DATA <= x"f656";
            when "00" & x"6d9" => DATA <= x"2400";
            when "00" & x"6da" => DATA <= x"6100";
            when "00" & x"6db" => DATA <= x"f61a";
            when "00" & x"6dc" => DATA <= x"2200";
            when "00" & x"6dd" => DATA <= x"6000";
            when "00" & x"6de" => DATA <= x"fc6a";
            when "00" & x"6df" => DATA <= x"2f00";
            when "00" & x"6e0" => DATA <= x"103c";
            when "00" & x"6e1" => DATA <= x"0012";
            when "00" & x"6e2" => DATA <= x"6100";
            when "00" & x"6e3" => DATA <= x"f61c";
            when "00" & x"6e4" => DATA <= x"201f";
            when "00" & x"6e5" => DATA <= x"6100";
            when "00" & x"6e6" => DATA <= x"f616";
            when "00" & x"6e7" => DATA <= x"4a40";
            when "00" & x"6e8" => DATA <= x"6600";
            when "00" & x"6e9" => DATA <= x"0012";
            when "00" & x"6ea" => DATA <= x"2f00";
            when "00" & x"6eb" => DATA <= x"1001";
            when "00" & x"6ec" => DATA <= x"6100";
            when "00" & x"6ed" => DATA <= x"f608";
            when "00" & x"6ee" => DATA <= x"6100";
            when "00" & x"6ef" => DATA <= x"f5f2";
            when "00" & x"6f0" => DATA <= x"201f";
            when "00" & x"6f1" => DATA <= x"4e75";
            when "00" & x"6f2" => DATA <= x"6100";
            when "00" & x"6f3" => DATA <= x"f650";
            when "00" & x"6f4" => DATA <= x"6000";
            when "00" & x"6f5" => DATA <= x"f5e6";
            when "00" & x"6f6" => DATA <= x"2800";
            when "00" & x"6f7" => DATA <= x"c8bc";
            when "00" & x"6f8" => DATA <= x"d000";
            when "00" & x"6f9" => DATA <= x"0000";
            when "00" & x"6fa" => DATA <= x"6000";
            when "00" & x"6fb" => DATA <= x"06f6";
            when "00" & x"6fc" => DATA <= x"2f05";
            when "00" & x"6fd" => DATA <= x"2f04";
            when "00" & x"6fe" => DATA <= x"2f01";
            when "00" & x"6ff" => DATA <= x"2f00";
            when "00" & x"700" => DATA <= x"2203";
            when "00" & x"701" => DATA <= x"700a";
            when "00" & x"702" => DATA <= x"6100";
            when "00" & x"703" => DATA <= x"04fa";
            when "00" & x"704" => DATA <= x"2801";
            when "00" & x"705" => DATA <= x"2202";
            when "00" & x"706" => DATA <= x"7009";
            when "00" & x"707" => DATA <= x"6100";
            when "00" & x"708" => DATA <= x"04f0";
            when "00" & x"709" => DATA <= x"2a01";
            when "00" & x"70a" => DATA <= x"221f";
            when "00" & x"70b" => DATA <= x"261f";
            when "00" & x"70c" => DATA <= x"7006";
            when "00" & x"70d" => DATA <= x"6100";
            when "00" & x"70e" => DATA <= x"04e4";
            when "00" & x"70f" => DATA <= x"2001";
            when "00" & x"710" => DATA <= x"2203";
            when "00" & x"711" => DATA <= x"2604";
            when "00" & x"712" => DATA <= x"2405";
            when "00" & x"713" => DATA <= x"281f";
            when "00" & x"714" => DATA <= x"2a1f";
            when "00" & x"715" => DATA <= x"023c";
            when "00" & x"716" => DATA <= x"00fd";
            when "00" & x"717" => DATA <= x"4e75";
            when "00" & x"718" => DATA <= x"203c";
            when "00" & x"719" => DATA <= x"0000";
            when "00" & x"71a" => DATA <= x"0600";
            when "00" & x"71b" => DATA <= x"223c";
            when "00" & x"71c" => DATA <= x"0000";
            when "00" & x"71d" => DATA <= x"0500";
            when "00" & x"71e" => DATA <= x"243c";
            when "00" & x"71f" => DATA <= x"0000";
            when "00" & x"720" => DATA <= x"052d";
            when "00" & x"721" => DATA <= x"4e75";
            when "00" & x"722" => DATA <= x"2f38";
            when "00" & x"723" => DATA <= x"04d0";
            when "00" & x"724" => DATA <= x"4e75";
            when "00" & x"725" => DATA <= x"2f03";
            when "00" & x"726" => DATA <= x"2f02";
            when "00" & x"727" => DATA <= x"2f01";
            when "00" & x"728" => DATA <= x"2f00";
            when "00" & x"729" => DATA <= x"2207";
            when "00" & x"72a" => DATA <= x"7004";
            when "00" & x"72b" => DATA <= x"6100";
            when "00" & x"72c" => DATA <= x"04a8";
            when "00" & x"72d" => DATA <= x"2e01";
            when "00" & x"72e" => DATA <= x"2206";
            when "00" & x"72f" => DATA <= x"7003";
            when "00" & x"730" => DATA <= x"6100";
            when "00" & x"731" => DATA <= x"049e";
            when "00" & x"732" => DATA <= x"2c01";
            when "00" & x"733" => DATA <= x"2205";
            when "00" & x"734" => DATA <= x"7002";
            when "00" & x"735" => DATA <= x"6100";
            when "00" & x"736" => DATA <= x"0494";
            when "00" & x"737" => DATA <= x"2a01";
            when "00" & x"738" => DATA <= x"2204";
            when "00" & x"739" => DATA <= x"7001";
            when "00" & x"73a" => DATA <= x"6100";
            when "00" & x"73b" => DATA <= x"048a";
            when "00" & x"73c" => DATA <= x"2801";
            when "00" & x"73d" => DATA <= x"221f";
            when "00" & x"73e" => DATA <= x"700b";
            when "00" & x"73f" => DATA <= x"6100";
            when "00" & x"740" => DATA <= x"0480";
            when "00" & x"741" => DATA <= x"2001";
            when "00" & x"742" => DATA <= x"221f";
            when "00" & x"743" => DATA <= x"2f00";
            when "00" & x"744" => DATA <= x"7000";
            when "00" & x"745" => DATA <= x"6100";
            when "00" & x"746" => DATA <= x"0474";
            when "00" & x"747" => DATA <= x"201f";
            when "00" & x"748" => DATA <= x"241f";
            when "00" & x"749" => DATA <= x"261f";
            when "00" & x"74a" => DATA <= x"023c";
            when "00" & x"74b" => DATA <= x"00fd";
            when "00" & x"74c" => DATA <= x"4e75";
            when "00" & x"74d" => DATA <= x"007c";
            when "00" & x"74e" => DATA <= x"0700";
            when "00" & x"74f" => DATA <= x"4e75";
            when "00" & x"750" => DATA <= x"027c";
            when "00" & x"751" => DATA <= x"f8ff";
            when "00" & x"752" => DATA <= x"4e75";
            when "00" & x"753" => DATA <= x"2f03";
            when "00" & x"754" => DATA <= x"2f02";
            when "00" & x"755" => DATA <= x"4282";
            when "00" & x"756" => DATA <= x"c343";
            when "00" & x"757" => DATA <= x"2200";
            when "00" & x"758" => DATA <= x"103c";
            when "00" & x"759" => DATA <= x"0007";
            when "00" & x"75a" => DATA <= x"6100";
            when "00" & x"75b" => DATA <= x"044a";
            when "00" & x"75c" => DATA <= x"c340";
            when "00" & x"75d" => DATA <= x"c741";
            when "00" & x"75e" => DATA <= x"241f";
            when "00" & x"75f" => DATA <= x"261f";
            when "00" & x"760" => DATA <= x"023c";
            when "00" & x"761" => DATA <= x"00fd";
            when "00" & x"762" => DATA <= x"4e75";
            when "00" & x"763" => DATA <= x"007c";
            when "00" & x"764" => DATA <= x"2000";
            when "00" & x"765" => DATA <= x"4e75";
            when "00" & x"766" => DATA <= x"2f03";
            when "00" & x"767" => DATA <= x"2f02";
            when "00" & x"768" => DATA <= x"4282";
            when "00" & x"769" => DATA <= x"c343";
            when "00" & x"76a" => DATA <= x"2200";
            when "00" & x"76b" => DATA <= x"103c";
            when "00" & x"76c" => DATA <= x"0008";
            when "00" & x"76d" => DATA <= x"6100";
            when "00" & x"76e" => DATA <= x"0424";
            when "00" & x"76f" => DATA <= x"c340";
            when "00" & x"770" => DATA <= x"c741";
            when "00" & x"771" => DATA <= x"241f";
            when "00" & x"772" => DATA <= x"261f";
            when "00" & x"773" => DATA <= x"023c";
            when "00" & x"774" => DATA <= x"00fd";
            when "00" & x"775" => DATA <= x"4e75";
            when "00" & x"776" => DATA <= x"2f03";
            when "00" & x"777" => DATA <= x"2f02";
            when "00" & x"778" => DATA <= x"2f01";
            when "00" & x"779" => DATA <= x"2200";
            when "00" & x"77a" => DATA <= x"103c";
            when "00" & x"77b" => DATA <= x"000c";
            when "00" & x"77c" => DATA <= x"6100";
            when "00" & x"77d" => DATA <= x"0406";
            when "00" & x"77e" => DATA <= x"2001";
            when "00" & x"77f" => DATA <= x"221f";
            when "00" & x"780" => DATA <= x"241f";
            when "00" & x"781" => DATA <= x"261f";
            when "00" & x"782" => DATA <= x"023c";
            when "00" & x"783" => DATA <= x"00fd";
            when "00" & x"784" => DATA <= x"4e75";
            when "00" & x"785" => DATA <= x"6100";
            when "00" & x"786" => DATA <= x"03fa";
            when "00" & x"787" => DATA <= x"2600";
            when "00" & x"788" => DATA <= x"7040";
            when "00" & x"789" => DATA <= x"2238";
            when "00" & x"78a" => DATA <= x"0600";
            when "00" & x"78b" => DATA <= x"6100";
            when "00" & x"78c" => DATA <= x"fccc";
            when "00" & x"78d" => DATA <= x"4280";
            when "00" & x"78e" => DATA <= x"4281";
            when "00" & x"78f" => DATA <= x"3038";
            when "00" & x"790" => DATA <= x"0600";
            when "00" & x"791" => DATA <= x"3238";
            when "00" & x"792" => DATA <= x"0600";
            when "00" & x"793" => DATA <= x"0480";
            when "00" & x"794" => DATA <= x"0000";
            when "00" & x"795" => DATA <= x"0280";
            when "00" & x"796" => DATA <= x"0481";
            when "00" & x"797" => DATA <= x"0000";
            when "00" & x"798" => DATA <= x"0200";
            when "00" & x"799" => DATA <= x"c1fc";
            when "00" & x"79a" => DATA <= x"0033";
            when "00" & x"79b" => DATA <= x"ed89";
            when "00" & x"79c" => DATA <= x"4282";
            when "00" & x"79d" => DATA <= x"0838";
            when "00" & x"79e" => DATA <= x"0007";
            when "00" & x"79f" => DATA <= x"0606";
            when "00" & x"7a0" => DATA <= x"6700";
            when "00" & x"7a1" => DATA <= x"0006";
            when "00" & x"7a2" => DATA <= x"08c2";
            when "00" & x"7a3" => DATA <= x"0000";
            when "00" & x"7a4" => DATA <= x"0838";
            when "00" & x"7a5" => DATA <= x"0006";
            when "00" & x"7a6" => DATA <= x"0606";
            when "00" & x"7a7" => DATA <= x"6700";
            when "00" & x"7a8" => DATA <= x"0006";
            when "00" & x"7a9" => DATA <= x"08c2";
            when "00" & x"7aa" => DATA <= x"0001";
            when "00" & x"7ab" => DATA <= x"0838";
            when "00" & x"7ac" => DATA <= x"0005";
            when "00" & x"7ad" => DATA <= x"0606";
            when "00" & x"7ae" => DATA <= x"6700";
            when "00" & x"7af" => DATA <= x"0006";
            when "00" & x"7b0" => DATA <= x"08c2";
            when "00" & x"7b1" => DATA <= x"0002";
            when "00" & x"7b2" => DATA <= x"023c";
            when "00" & x"7b3" => DATA <= x"00fd";
            when "00" & x"7b4" => DATA <= x"4e75";
            when "00" & x"7b5" => DATA <= x"103c";
            when "00" & x"7b6" => DATA <= x"0080";
            when "00" & x"7b7" => DATA <= x"123c";
            when "00" & x"7b8" => DATA <= x"0007";
            when "00" & x"7b9" => DATA <= x"143c";
            when "00" & x"7ba" => DATA <= x"0000";
            when "00" & x"7bb" => DATA <= x"6100";
            when "00" & x"7bc" => DATA <= x"fb5a";
            when "00" & x"7bd" => DATA <= x"103c";
            when "00" & x"7be" => DATA <= x"0080";
            when "00" & x"7bf" => DATA <= x"123c";
            when "00" & x"7c0" => DATA <= x"0008";
            when "00" & x"7c1" => DATA <= x"143c";
            when "00" & x"7c2" => DATA <= x"0000";
            when "00" & x"7c3" => DATA <= x"6100";
            when "00" & x"7c4" => DATA <= x"fb4a";
            when "00" & x"7c5" => DATA <= x"103c";
            when "00" & x"7c6" => DATA <= x"0080";
            when "00" & x"7c7" => DATA <= x"123c";
            when "00" & x"7c8" => DATA <= x"0009";
            when "00" & x"7c9" => DATA <= x"143c";
            when "00" & x"7ca" => DATA <= x"0000";
            when "00" & x"7cb" => DATA <= x"6100";
            when "00" & x"7cc" => DATA <= x"fb3a";
            when "00" & x"7cd" => DATA <= x"103c";
            when "00" & x"7ce" => DATA <= x"0081";
            when "00" & x"7cf" => DATA <= x"123c";
            when "00" & x"7d0" => DATA <= x"00f6";
            when "00" & x"7d1" => DATA <= x"143c";
            when "00" & x"7d2" => DATA <= x"00ff";
            when "00" & x"7d3" => DATA <= x"6100";
            when "00" & x"7d4" => DATA <= x"fb2a";
            when "00" & x"7d5" => DATA <= x"103c";
            when "00" & x"7d6" => DATA <= x"0081";
            when "00" & x"7d7" => DATA <= x"123c";
            when "00" & x"7d8" => DATA <= x"00f5";
            when "00" & x"7d9" => DATA <= x"143c";
            when "00" & x"7da" => DATA <= x"00ff";
            when "00" & x"7db" => DATA <= x"6100";
            when "00" & x"7dc" => DATA <= x"fb1a";
            when "00" & x"7dd" => DATA <= x"103c";
            when "00" & x"7de" => DATA <= x"0081";
            when "00" & x"7df" => DATA <= x"123c";
            when "00" & x"7e0" => DATA <= x"00f4";
            when "00" & x"7e1" => DATA <= x"143c";
            when "00" & x"7e2" => DATA <= x"00ff";
            when "00" & x"7e3" => DATA <= x"6100";
            when "00" & x"7e4" => DATA <= x"fb0a";
            when "00" & x"7e5" => DATA <= x"4e75";
            when "00" & x"7e6" => DATA <= x"2f0e";
            when "00" & x"7e7" => DATA <= x"2f07";
            when "00" & x"7e8" => DATA <= x"2f06";
            when "00" & x"7e9" => DATA <= x"2f04";
            when "00" & x"7ea" => DATA <= x"2f03";
            when "00" & x"7eb" => DATA <= x"2f00";
            when "00" & x"7ec" => DATA <= x"7eff";
            when "00" & x"7ed" => DATA <= x"0800";
            when "00" & x"7ee" => DATA <= x"001d";
            when "00" & x"7ef" => DATA <= x"6700";
            when "00" & x"7f0" => DATA <= x"0004";
            when "00" & x"7f1" => DATA <= x"2e02";
            when "00" & x"7f2" => DATA <= x"0280";
            when "00" & x"7f3" => DATA <= x"0000";
            when "00" & x"7f4" => DATA <= x"00ff";
            when "00" & x"7f5" => DATA <= x"4a80";
            when "00" & x"7f6" => DATA <= x"6600";
            when "00" & x"7f7" => DATA <= x"0004";
            when "00" & x"7f8" => DATA <= x"700a";
            when "00" & x"7f9" => DATA <= x"b0bc";
            when "00" & x"7fa" => DATA <= x"0000";
            when "00" & x"7fb" => DATA <= x"0002";
            when "00" & x"7fc" => DATA <= x"6500";
            when "00" & x"7fd" => DATA <= x"00a0";
            when "00" & x"7fe" => DATA <= x"b0bc";
            when "00" & x"7ff" => DATA <= x"0000";
            when "00" & x"800" => DATA <= x"0024";
            when "00" & x"801" => DATA <= x"6200";
            when "00" & x"802" => DATA <= x"0096";
            when "00" & x"803" => DATA <= x"2c00";
            when "00" & x"804" => DATA <= x"4282";
            when "00" & x"805" => DATA <= x"2c41";
            when "00" & x"806" => DATA <= x"6100";
            when "00" & x"807" => DATA <= x"1712";
            when "00" & x"808" => DATA <= x"528e";
            when "00" & x"809" => DATA <= x"b03c";
            when "00" & x"80a" => DATA <= x"0026";
            when "00" & x"80b" => DATA <= x"6600";
            when "00" & x"80c" => DATA <= x"000a";
            when "00" & x"80d" => DATA <= x"7c10";
            when "00" & x"80e" => DATA <= x"528e";
            when "00" & x"80f" => DATA <= x"6000";
            when "00" & x"810" => DATA <= x"000e";
            when "00" & x"811" => DATA <= x"b03c";
            when "00" & x"812" => DATA <= x"0024";
            when "00" & x"813" => DATA <= x"6600";
            when "00" & x"814" => DATA <= x"0006";
            when "00" & x"815" => DATA <= x"7c10";
            when "00" & x"816" => DATA <= x"528e";
            when "00" & x"817" => DATA <= x"0c00";
            when "00" & x"818" => DATA <= x"0039";
            when "00" & x"819" => DATA <= x"6300";
            when "00" & x"81a" => DATA <= x"0008";
            when "00" & x"81b" => DATA <= x"0200";
            when "00" & x"81c" => DATA <= x"00df";
            when "00" & x"81d" => DATA <= x"5f00";
            when "00" & x"81e" => DATA <= x"0400";
            when "00" & x"81f" => DATA <= x"0030";
            when "00" & x"820" => DATA <= x"6b00";
            when "00" & x"821" => DATA <= x"0030";
            when "00" & x"822" => DATA <= x"b006";
            when "00" & x"823" => DATA <= x"6200";
            when "00" & x"824" => DATA <= x"002a";
            when "00" & x"825" => DATA <= x"bcbc";
            when "00" & x"826" => DATA <= x"0000";
            when "00" & x"827" => DATA <= x"0010";
            when "00" & x"828" => DATA <= x"6600";
            when "00" & x"829" => DATA <= x"000a";
            when "00" & x"82a" => DATA <= x"e98a";
            when "00" & x"82b" => DATA <= x"d480";
            when "00" & x"82c" => DATA <= x"101e";
            when "00" & x"82d" => DATA <= x"60d2";
            when "00" & x"82e" => DATA <= x"2606";
            when "00" & x"82f" => DATA <= x"5583";
            when "00" & x"830" => DATA <= x"2802";
            when "00" & x"831" => DATA <= x"d484";
            when "00" & x"832" => DATA <= x"6500";
            when "00" & x"833" => DATA <= x"0048";
            when "00" & x"834" => DATA <= x"51cb";
            when "00" & x"835" => DATA <= x"fff8";
            when "00" & x"836" => DATA <= x"d480";
            when "00" & x"837" => DATA <= x"101e";
            when "00" & x"838" => DATA <= x"60bc";
            when "00" & x"839" => DATA <= x"4a82";
            when "00" & x"83a" => DATA <= x"6700";
            when "00" & x"83b" => DATA <= x"002e";
            when "00" & x"83c" => DATA <= x"4a87";
            when "00" & x"83d" => DATA <= x"6700";
            when "00" & x"83e" => DATA <= x"0008";
            when "00" & x"83f" => DATA <= x"b087";
            when "00" & x"840" => DATA <= x"6200";
            when "00" & x"841" => DATA <= x"002c";
            when "00" & x"842" => DATA <= x"220e";
            when "00" & x"843" => DATA <= x"5381";
            when "00" & x"844" => DATA <= x"201f";
            when "00" & x"845" => DATA <= x"261f";
            when "00" & x"846" => DATA <= x"281f";
            when "00" & x"847" => DATA <= x"2c1f";
            when "00" & x"848" => DATA <= x"2e1f";
            when "00" & x"849" => DATA <= x"2c5f";
            when "00" & x"84a" => DATA <= x"023c";
            when "00" & x"84b" => DATA <= x"00fd";
            when "00" & x"84c" => DATA <= x"4e75";
            when "00" & x"84d" => DATA <= x"203c";
            when "00" & x"84e" => DATA <= x"003f";
            when "00" & x"84f" => DATA <= x"2de8";
            when "00" & x"850" => DATA <= x"6000";
            when "00" & x"851" => DATA <= x"0012";
            when "00" & x"852" => DATA <= x"203c";
            when "00" & x"853" => DATA <= x"003f";
            when "00" & x"854" => DATA <= x"2df8";
            when "00" & x"855" => DATA <= x"6000";
            when "00" & x"856" => DATA <= x"0008";
            when "00" & x"857" => DATA <= x"203c";
            when "00" & x"858" => DATA <= x"003f";
            when "00" & x"859" => DATA <= x"2e08";
            when "00" & x"85a" => DATA <= x"261f";
            when "00" & x"85b" => DATA <= x"261f";
            when "00" & x"85c" => DATA <= x"281f";
            when "00" & x"85d" => DATA <= x"2c1f";
            when "00" & x"85e" => DATA <= x"2e1f";
            when "00" & x"85f" => DATA <= x"2c5f";
            when "00" & x"860" => DATA <= x"003c";
            when "00" & x"861" => DATA <= x"0002";
            when "00" & x"862" => DATA <= x"4e75";
            when "00" & x"863" => DATA <= x"2f00";
            when "00" & x"864" => DATA <= x"2f01";
            when "00" & x"865" => DATA <= x"6100";
            when "00" & x"866" => DATA <= x"07bc";
            when "00" & x"867" => DATA <= x"2401";
            when "00" & x"868" => DATA <= x"221f";
            when "00" & x"869" => DATA <= x"201f";
            when "00" & x"86a" => DATA <= x"4e75";
            when "00" & x"86b" => DATA <= x"b03c";
            when "00" & x"86c" => DATA <= x"003a";
            when "00" & x"86d" => DATA <= x"6200";
            when "00" & x"86e" => DATA <= x"001c";
            when "00" & x"86f" => DATA <= x"2f0e";
            when "00" & x"870" => DATA <= x"d040";
            when "00" & x"871" => DATA <= x"d040";
            when "00" & x"872" => DATA <= x"2c79";
            when "00" & x"873" => DATA <= x"003f";
            when "00" & x"874" => DATA <= x"36f8";
            when "00" & x"875" => DATA <= x"ddc0";
            when "00" & x"876" => DATA <= x"4dd6";
            when "00" & x"877" => DATA <= x"4e96";
            when "00" & x"878" => DATA <= x"2c5f";
            when "00" & x"879" => DATA <= x"023c";
            when "00" & x"87a" => DATA <= x"00fd";
            when "00" & x"87b" => DATA <= x"4e75";
            when "00" & x"87c" => DATA <= x"203c";
            when "00" & x"87d" => DATA <= x"003f";
            when "00" & x"87e" => DATA <= x"2ef4";
            when "00" & x"87f" => DATA <= x"003c";
            when "00" & x"880" => DATA <= x"0002";
            when "00" & x"881" => DATA <= x"4e75";
            when "00" & x"882" => DATA <= x"103c";
            when "00" & x"883" => DATA <= x"008b";
            when "00" & x"884" => DATA <= x"6100";
            when "00" & x"885" => DATA <= x"f9c8";
            when "00" & x"886" => DATA <= x"103c";
            when "00" & x"887" => DATA <= x"0010";
            when "00" & x"888" => DATA <= x"4e75";
            when "00" & x"889" => DATA <= x"7000";
            when "00" & x"88a" => DATA <= x"7200";
            when "00" & x"88b" => DATA <= x"6100";
            when "00" & x"88c" => DATA <= x"fbb2";
            when "00" & x"88d" => DATA <= x"103c";
            when "00" & x"88e" => DATA <= x"0016";
            when "00" & x"88f" => DATA <= x"4e75";
            when "00" & x"890" => DATA <= x"2f38";
            when "00" & x"891" => DATA <= x"0404";
            when "00" & x"892" => DATA <= x"4e75";
            when "00" & x"893" => DATA <= x"0838";
            when "00" & x"894" => DATA <= x"0006";
            when "00" & x"895" => DATA <= x"0535";
            when "00" & x"896" => DATA <= x"6600";
            when "00" & x"897" => DATA <= x"0008";
            when "00" & x"898" => DATA <= x"023c";
            when "00" & x"899" => DATA <= x"00fe";
            when "00" & x"89a" => DATA <= x"4e75";
            when "00" & x"89b" => DATA <= x"003c";
            when "00" & x"89c" => DATA <= x"0001";
            when "00" & x"89d" => DATA <= x"4e75";
            when "00" & x"89e" => DATA <= x"2f04";
            when "00" & x"89f" => DATA <= x"7801";
            when "00" & x"8a0" => DATA <= x"2f0e";
            when "00" & x"8a1" => DATA <= x"2c79";
            when "00" & x"8a2" => DATA <= x"0000";
            when "00" & x"8a3" => DATA <= x"048c";
            when "00" & x"8a4" => DATA <= x"4e96";
            when "00" & x"8a5" => DATA <= x"2c5f";
            when "00" & x"8a6" => DATA <= x"281f";
            when "00" & x"8a7" => DATA <= x"4e75";
            when "00" & x"8a8" => DATA <= x"4e75";
            when "00" & x"8a9" => DATA <= x"b0bc";
            when "00" & x"8aa" => DATA <= x"0000";
            when "00" & x"8ab" => DATA <= x"04ff";
            when "00" & x"8ac" => DATA <= x"6200";
            when "00" & x"8ad" => DATA <= x"0040";
            when "00" & x"8ae" => DATA <= x"b2bc";
            when "00" & x"8af" => DATA <= x"0000";
            when "00" & x"8b0" => DATA <= x"03ff";
            when "00" & x"8b1" => DATA <= x"6200";
            when "00" & x"8b2" => DATA <= x"0036";
            when "00" & x"8b3" => DATA <= x"2f00";
            when "00" & x"8b4" => DATA <= x"2f01";
            when "00" & x"8b5" => DATA <= x"31c0";
            when "00" & x"8b6" => DATA <= x"0600";
            when "00" & x"8b7" => DATA <= x"31c1";
            when "00" & x"8b8" => DATA <= x"0602";
            when "00" & x"8b9" => DATA <= x"223c";
            when "00" & x"8ba" => DATA <= x"0000";
            when "00" & x"8bb" => DATA <= x"0600";
            when "00" & x"8bc" => DATA <= x"7009";
            when "00" & x"8bd" => DATA <= x"6100";
            when "00" & x"8be" => DATA <= x"fa68";
            when "00" & x"8bf" => DATA <= x"7400";
            when "00" & x"8c0" => DATA <= x"7600";
            when "00" & x"8c1" => DATA <= x"1438";
            when "00" & x"8c2" => DATA <= x"0604";
            when "00" & x"8c3" => DATA <= x"221f";
            when "00" & x"8c4" => DATA <= x"201f";
            when "00" & x"8c5" => DATA <= x"b43c";
            when "00" & x"8c6" => DATA <= x"00ff";
            when "00" & x"8c7" => DATA <= x"6700";
            when "00" & x"8c8" => DATA <= x"000a";
            when "00" & x"8c9" => DATA <= x"7800";
            when "00" & x"8ca" => DATA <= x"023c";
            when "00" & x"8cb" => DATA <= x"00fd";
            when "00" & x"8cc" => DATA <= x"4e75";
            when "00" & x"8cd" => DATA <= x"203c";
            when "00" & x"8ce" => DATA <= x"003f";
            when "00" & x"8cf" => DATA <= x"2d64";
            when "00" & x"8d0" => DATA <= x"78ff";
            when "00" & x"8d1" => DATA <= x"003c";
            when "00" & x"8d2" => DATA <= x"0002";
            when "00" & x"8d3" => DATA <= x"4e75";
            when "00" & x"8d4" => DATA <= x"b5fc";
            when "00" & x"8d5" => DATA <= x"0000";
            when "00" & x"8d6" => DATA <= x"002f";
            when "00" & x"8d7" => DATA <= x"6200";
            when "00" & x"8d8" => DATA <= x"0018";
            when "00" & x"8d9" => DATA <= x"2f0a";
            when "00" & x"8da" => DATA <= x"d4ca";
            when "00" & x"8db" => DATA <= x"d4ca";
            when "00" & x"8dc" => DATA <= x"d5f8";
            when "00" & x"8dd" => DATA <= x"0000";
            when "00" & x"8de" => DATA <= x"45d2";
            when "00" & x"8df" => DATA <= x"4e92";
            when "00" & x"8e0" => DATA <= x"245f";
            when "00" & x"8e1" => DATA <= x"023c";
            when "00" & x"8e2" => DATA <= x"00fd";
            when "00" & x"8e3" => DATA <= x"4e75";
            when "00" & x"8e4" => DATA <= x"203c";
            when "00" & x"8e5" => DATA <= x"003f";
            when "00" & x"8e6" => DATA <= x"2e48";
            when "00" & x"8e7" => DATA <= x"003c";
            when "00" & x"8e8" => DATA <= x"0002";
            when "00" & x"8e9" => DATA <= x"4e75";
            when "00" & x"8ea" => DATA <= x"2f00";
            when "00" & x"8eb" => DATA <= x"2f01";
            when "00" & x"8ec" => DATA <= x"203c";
            when "00" & x"8ed" => DATA <= x"003f";
            when "00" & x"8ee" => DATA <= x"2822";
            when "00" & x"8ef" => DATA <= x"720b";
            when "00" & x"8f0" => DATA <= x"6100";
            when "00" & x"8f1" => DATA <= x"018c";
            when "00" & x"8f2" => DATA <= x"221f";
            when "00" & x"8f3" => DATA <= x"201f";
            when "00" & x"8f4" => DATA <= x"023c";
            when "00" & x"8f5" => DATA <= x"00fd";
            when "00" & x"8f6" => DATA <= x"4e75";
            when "00" & x"8f7" => DATA <= x"2f00";
            when "00" & x"8f8" => DATA <= x"2f01";
            when "00" & x"8f9" => DATA <= x"203c";
            when "00" & x"8fa" => DATA <= x"003f";
            when "00" & x"8fb" => DATA <= x"282d";
            when "00" & x"8fc" => DATA <= x"720b";
            when "00" & x"8fd" => DATA <= x"6100";
            when "00" & x"8fe" => DATA <= x"0172";
            when "00" & x"8ff" => DATA <= x"221f";
            when "00" & x"900" => DATA <= x"201f";
            when "00" & x"901" => DATA <= x"023c";
            when "00" & x"902" => DATA <= x"00fd";
            when "00" & x"903" => DATA <= x"4e75";
            when "00" & x"904" => DATA <= x"2f0e";
            when "00" & x"905" => DATA <= x"2f09";
            when "00" & x"906" => DATA <= x"2f01";
            when "00" & x"907" => DATA <= x"2f00";
            when "00" & x"908" => DATA <= x"2c41";
            when "00" & x"909" => DATA <= x"0280";
            when "00" & x"90a" => DATA <= x"0002";
            when "00" & x"90b" => DATA <= x"0000";
            when "00" & x"90c" => DATA <= x"6700";
            when "00" & x"90d" => DATA <= x"000c";
            when "00" & x"90e" => DATA <= x"5382";
            when "00" & x"90f" => DATA <= x"6b00";
            when "00" & x"910" => DATA <= x"005c";
            when "00" & x"911" => DATA <= x"1cfc";
            when "00" & x"912" => DATA <= x"0058";
            when "00" & x"913" => DATA <= x"43f9";
            when "00" & x"914" => DATA <= x"003f";
            when "00" & x"915" => DATA <= x"2f50";
            when "00" & x"916" => DATA <= x"b099";
            when "00" & x"917" => DATA <= x"6700";
            when "00" & x"918" => DATA <= x"0014";
            when "00" & x"919" => DATA <= x"2219";
            when "00" & x"91a" => DATA <= x"b23c";
            when "00" & x"91b" => DATA <= x"00ff";
            when "00" & x"91c" => DATA <= x"6700";
            when "00" & x"91d" => DATA <= x"0020";
            when "00" & x"91e" => DATA <= x"b23c";
            when "00" & x"91f" => DATA <= x"0000";
            when "00" & x"920" => DATA <= x"66f0";
            when "00" & x"921" => DATA <= x"60e8";
            when "00" & x"922" => DATA <= x"2019";
            when "00" & x"923" => DATA <= x"5382";
            when "00" & x"924" => DATA <= x"6b00";
            when "00" & x"925" => DATA <= x"0032";
            when "00" & x"926" => DATA <= x"1cd9";
            when "00" & x"927" => DATA <= x"66f6";
            when "00" & x"928" => DATA <= x"201f";
            when "00" & x"929" => DATA <= x"221f";
            when "00" & x"92a" => DATA <= x"225f";
            when "00" & x"92b" => DATA <= x"2c5f";
            when "00" & x"92c" => DATA <= x"4e75";
            when "00" & x"92d" => DATA <= x"0c81";
            when "00" & x"92e" => DATA <= x"0000";
            when "00" & x"92f" => DATA <= x"000d";
            when "00" & x"930" => DATA <= x"6500";
            when "00" & x"931" => DATA <= x"001a";
            when "00" & x"932" => DATA <= x"2cfc";
            when "00" & x"933" => DATA <= x"4f53";
            when "00" & x"934" => DATA <= x"5f55";
            when "00" & x"935" => DATA <= x"2cfc";
            when "00" & x"936" => DATA <= x"6e64";
            when "00" & x"937" => DATA <= x"6566";
            when "00" & x"938" => DATA <= x"2cfc";
            when "00" & x"939" => DATA <= x"696e";
            when "00" & x"93a" => DATA <= x"6564";
            when "00" & x"93b" => DATA <= x"1cfc";
            when "00" & x"93c" => DATA <= x"0000";
            when "00" & x"93d" => DATA <= x"60d4";
            when "00" & x"93e" => DATA <= x"003c";
            when "00" & x"93f" => DATA <= x"0002";
            when "00" & x"940" => DATA <= x"2ebc";
            when "00" & x"941" => DATA <= x"003f";
            when "00" & x"942" => DATA <= x"2e80";
            when "00" & x"943" => DATA <= x"60c8";
            when "00" & x"944" => DATA <= x"2f0e";
            when "00" & x"945" => DATA <= x"2f0d";
            when "00" & x"946" => DATA <= x"2f01";
            when "00" & x"947" => DATA <= x"4bf9";
            when "00" & x"948" => DATA <= x"003f";
            when "00" & x"949" => DATA <= x"2f50";
            when "00" & x"94a" => DATA <= x"2c57";
            when "00" & x"94b" => DATA <= x"201d";
            when "00" & x"94c" => DATA <= x"588d";
            when "00" & x"94d" => DATA <= x"bd8d";
            when "00" & x"94e" => DATA <= x"6600";
            when "00" & x"94f" => DATA <= x"0010";
            when "00" & x"950" => DATA <= x"4a2d";
            when "00" & x"951" => DATA <= x"ffff";
            when "00" & x"952" => DATA <= x"66f4";
            when "00" & x"953" => DATA <= x"221f";
            when "00" & x"954" => DATA <= x"2a5f";
            when "00" & x"955" => DATA <= x"2c5f";
            when "00" & x"956" => DATA <= x"4e75";
            when "00" & x"957" => DATA <= x"201d";
            when "00" & x"958" => DATA <= x"4a00";
            when "00" & x"959" => DATA <= x"66fa";
            when "00" & x"95a" => DATA <= x"b03c";
            when "00" & x"95b" => DATA <= x"00ff";
            when "00" & x"95c" => DATA <= x"66da";
            when "00" & x"95d" => DATA <= x"221f";
            when "00" & x"95e" => DATA <= x"2a5f";
            when "00" & x"95f" => DATA <= x"2c5f";
            when "00" & x"960" => DATA <= x"203c";
            when "00" & x"961" => DATA <= x"003f";
            when "00" & x"962" => DATA <= x"2e94";
            when "00" & x"963" => DATA <= x"003c";
            when "00" & x"964" => DATA <= x"0002";
            when "00" & x"965" => DATA <= x"4e75";
            when "00" & x"966" => DATA <= x"4a80";
            when "00" & x"967" => DATA <= x"6d00";
            when "00" & x"968" => DATA <= x"0010";
            when "00" & x"969" => DATA <= x"b2b8";
            when "00" & x"96a" => DATA <= x"0508";
            when "00" & x"96b" => DATA <= x"6200";
            when "00" & x"96c" => DATA <= x"0008";
            when "00" & x"96d" => DATA <= x"023c";
            when "00" & x"96e" => DATA <= x"00fe";
            when "00" & x"96f" => DATA <= x"4e75";
            when "00" & x"970" => DATA <= x"003c";
            when "00" & x"971" => DATA <= x"0001";
            when "00" & x"972" => DATA <= x"4e75";
            when "00" & x"973" => DATA <= x"0c80";
            when "00" & x"974" => DATA <= x"0000";
            when "00" & x"975" => DATA <= x"0007";
            when "00" & x"976" => DATA <= x"6200";
            when "00" & x"977" => DATA <= x"0008";
            when "00" & x"978" => DATA <= x"023c";
            when "00" & x"979" => DATA <= x"00fe";
            when "00" & x"97a" => DATA <= x"4e75";
            when "00" & x"97b" => DATA <= x"70ff";
            when "00" & x"97c" => DATA <= x"72fe";
            when "00" & x"97d" => DATA <= x"003c";
            when "00" & x"97e" => DATA <= x"0001";
            when "00" & x"97f" => DATA <= x"4e75";
            when "00" & x"980" => DATA <= x"2f38";
            when "00" & x"981" => DATA <= x"0478";
            when "00" & x"982" => DATA <= x"4e75";
            when "00" & x"983" => DATA <= x"2f01";
            when "00" & x"984" => DATA <= x"7001";
            when "00" & x"985" => DATA <= x"223c";
            when "00" & x"986" => DATA <= x"0000";
            when "00" & x"987" => DATA <= x"0600";
            when "00" & x"988" => DATA <= x"6100";
            when "00" & x"989" => DATA <= x"f8d2";
            when "00" & x"98a" => DATA <= x"2038";
            when "00" & x"98b" => DATA <= x"0600";
            when "00" & x"98c" => DATA <= x"90b8";
            when "00" & x"98d" => DATA <= x"0528";
            when "00" & x"98e" => DATA <= x"221f";
            when "00" & x"98f" => DATA <= x"4e75";
            when "00" & x"990" => DATA <= x"b0bc";
            when "00" & x"991" => DATA <= x"0000";
            when "00" & x"992" => DATA <= x"04ff";
            when "00" & x"993" => DATA <= x"6200";
            when "00" & x"994" => DATA <= x"0038";
            when "00" & x"995" => DATA <= x"b2bc";
            when "00" & x"996" => DATA <= x"0000";
            when "00" & x"997" => DATA <= x"03ff";
            when "00" & x"998" => DATA <= x"6200";
            when "00" & x"999" => DATA <= x"002e";
            when "00" & x"99a" => DATA <= x"2f00";
            when "00" & x"99b" => DATA <= x"7019";
            when "00" & x"99c" => DATA <= x"6100";
            when "00" & x"99d" => DATA <= x"f6ac";
            when "00" & x"99e" => DATA <= x"201f";
            when "00" & x"99f" => DATA <= x"6100";
            when "00" & x"9a0" => DATA <= x"f6a6";
            when "00" & x"9a1" => DATA <= x"3001";
            when "00" & x"9a2" => DATA <= x"6100";
            when "00" & x"9a3" => DATA <= x"f6a0";
            when "00" & x"9a4" => DATA <= x"e088";
            when "00" & x"9a5" => DATA <= x"6100";
            when "00" & x"9a6" => DATA <= x"f69a";
            when "00" & x"9a7" => DATA <= x"3002";
            when "00" & x"9a8" => DATA <= x"6100";
            when "00" & x"9a9" => DATA <= x"f694";
            when "00" & x"9aa" => DATA <= x"e088";
            when "00" & x"9ab" => DATA <= x"6100";
            when "00" & x"9ac" => DATA <= x"f68e";
            when "00" & x"9ad" => DATA <= x"023c";
            when "00" & x"9ae" => DATA <= x"00fd";
            when "00" & x"9af" => DATA <= x"4e75";
            when "00" & x"9b0" => DATA <= x"203c";
            when "00" & x"9b1" => DATA <= x"003f";
            when "00" & x"9b2" => DATA <= x"2d64";
            when "00" & x"9b3" => DATA <= x"78ff";
            when "00" & x"9b4" => DATA <= x"003c";
            when "00" & x"9b5" => DATA <= x"0002";
            when "00" & x"9b6" => DATA <= x"4e75";
            when "00" & x"9b7" => DATA <= x"0c81";
            when "00" & x"9b8" => DATA <= x"0000";
            when "00" & x"9b9" => DATA <= x"0000";
            when "00" & x"9ba" => DATA <= x"6700";
            when "00" & x"9bb" => DATA <= x"001c";
            when "00" & x"9bc" => DATA <= x"5341";
            when "00" & x"9bd" => DATA <= x"2f08";
            when "00" & x"9be" => DATA <= x"2f00";
            when "00" & x"9bf" => DATA <= x"2f01";
            when "00" & x"9c0" => DATA <= x"2040";
            when "00" & x"9c1" => DATA <= x"1018";
            when "00" & x"9c2" => DATA <= x"6100";
            when "00" & x"9c3" => DATA <= x"f660";
            when "00" & x"9c4" => DATA <= x"51c9";
            when "00" & x"9c5" => DATA <= x"fff8";
            when "00" & x"9c6" => DATA <= x"221f";
            when "00" & x"9c7" => DATA <= x"201f";
            when "00" & x"9c8" => DATA <= x"205f";
            when "00" & x"9c9" => DATA <= x"4e75";
            when "00" & x"9ca" => DATA <= x"2f0e";
            when "00" & x"9cb" => DATA <= x"2f0d";
            when "00" & x"9cc" => DATA <= x"4a80";
            when "00" & x"9cd" => DATA <= x"6700";
            when "00" & x"9ce" => DATA <= x"000e";
            when "00" & x"9cf" => DATA <= x"2c40";
            when "00" & x"9d0" => DATA <= x"2a7c";
            when "00" & x"9d1" => DATA <= x"0000";
            when "00" & x"9d2" => DATA <= x"0600";
            when "00" & x"9d3" => DATA <= x"1ade";
            when "00" & x"9d4" => DATA <= x"66fc";
            when "00" & x"9d5" => DATA <= x"4a81";
            when "00" & x"9d6" => DATA <= x"6700";
            when "00" & x"9d7" => DATA <= x"0016";
            when "00" & x"9d8" => DATA <= x"2f02";
            when "00" & x"9d9" => DATA <= x"7404";
            when "00" & x"9da" => DATA <= x"2c41";
            when "00" & x"9db" => DATA <= x"2a7c";
            when "00" & x"9dc" => DATA <= x"0000";
            when "00" & x"9dd" => DATA <= x"052d";
            when "00" & x"9de" => DATA <= x"1ade";
            when "00" & x"9df" => DATA <= x"5382";
            when "00" & x"9e0" => DATA <= x"6afa";
            when "00" & x"9e1" => DATA <= x"241f";
            when "00" & x"9e2" => DATA <= x"2a5f";
            when "00" & x"9e3" => DATA <= x"2c5f";
            when "00" & x"9e4" => DATA <= x"4e75";
            when "00" & x"9e5" => DATA <= x"2f02";
            when "00" & x"9e6" => DATA <= x"2f01";
            when "00" & x"9e7" => DATA <= x"2f00";
            when "00" & x"9e8" => DATA <= x"2203";
            when "00" & x"9e9" => DATA <= x"7004";
            when "00" & x"9ea" => DATA <= x"6100";
            when "00" & x"9eb" => DATA <= x"fbf4";
            when "00" & x"9ec" => DATA <= x"201f";
            when "00" & x"9ed" => DATA <= x"221f";
            when "00" & x"9ee" => DATA <= x"241f";
            when "00" & x"9ef" => DATA <= x"6000";
            when "00" & x"9f0" => DATA <= x"fa64";
            when "00" & x"9f1" => DATA <= x"b07c";
            when "00" & x"9f2" => DATA <= x"0010";
            when "00" & x"9f3" => DATA <= x"6300";
            when "00" & x"9f4" => DATA <= x"000e";
            when "00" & x"9f5" => DATA <= x"203c";
            when "00" & x"9f6" => DATA <= x"003f";
            when "00" & x"9f7" => DATA <= x"2e1c";
            when "00" & x"9f8" => DATA <= x"003c";
            when "00" & x"9f9" => DATA <= x"0002";
            when "00" & x"9fa" => DATA <= x"4e75";
            when "00" & x"9fb" => DATA <= x"41f9";
            when "00" & x"9fc" => DATA <= x"003f";
            when "00" & x"9fd" => DATA <= x"362c";
            when "00" & x"9fe" => DATA <= x"e588";
            when "00" & x"9ff" => DATA <= x"d1c0";
            when "00" & x"a00" => DATA <= x"d1c0";
            when "00" & x"a01" => DATA <= x"d1c0";
            when "00" & x"a02" => DATA <= x"2218";
            when "00" & x"a03" => DATA <= x"6700";
            when "00" & x"a04" => DATA <= x"11ea";
            when "00" & x"a05" => DATA <= x"0681";
            when "00" & x"a06" => DATA <= x"003f";
            when "00" & x"a07" => DATA <= x"0000";
            when "00" & x"a08" => DATA <= x"2418";
            when "00" & x"a09" => DATA <= x"6700";
            when "00" & x"a0a" => DATA <= x"0008";
            when "00" & x"a0b" => DATA <= x"0682";
            when "00" & x"a0c" => DATA <= x"003f";
            when "00" & x"a0d" => DATA <= x"0000";
            when "00" & x"a0e" => DATA <= x"2618";
            when "00" & x"a0f" => DATA <= x"6700";
            when "00" & x"a10" => DATA <= x"0008";
            when "00" & x"a11" => DATA <= x"0683";
            when "00" & x"a12" => DATA <= x"003f";
            when "00" & x"a13" => DATA <= x"0000";
            when "00" & x"a14" => DATA <= x"4e75";
            when "00" & x"a15" => DATA <= x"b0bc";
            when "00" & x"a16" => DATA <= x"0000";
            when "00" & x"a17" => DATA <= x"04ff";
            when "00" & x"a18" => DATA <= x"6200";
            when "00" & x"a19" => DATA <= x"005c";
            when "00" & x"a1a" => DATA <= x"b2bc";
            when "00" & x"a1b" => DATA <= x"0000";
            when "00" & x"a1c" => DATA <= x"03ff";
            when "00" & x"a1d" => DATA <= x"6200";
            when "00" & x"a1e" => DATA <= x"0052";
            when "00" & x"a1f" => DATA <= x"2f00";
            when "00" & x"a20" => DATA <= x"2f01";
            when "00" & x"a21" => DATA <= x"103c";
            when "00" & x"a22" => DATA <= x"0017";
            when "00" & x"a23" => DATA <= x"6100";
            when "00" & x"a24" => DATA <= x"f59e";
            when "00" & x"a25" => DATA <= x"103c";
            when "00" & x"a26" => DATA <= x"0011";
            when "00" & x"a27" => DATA <= x"6100";
            when "00" & x"a28" => DATA <= x"f596";
            when "00" & x"a29" => DATA <= x"103c";
            when "00" & x"a2a" => DATA <= x"0006";
            when "00" & x"a2b" => DATA <= x"6100";
            when "00" & x"a2c" => DATA <= x"f58e";
            when "00" & x"a2d" => DATA <= x"201f";
            when "00" & x"a2e" => DATA <= x"e098";
            when "00" & x"a2f" => DATA <= x"6100";
            when "00" & x"a30" => DATA <= x"f586";
            when "00" & x"a31" => DATA <= x"e198";
            when "00" & x"a32" => DATA <= x"6100";
            when "00" & x"a33" => DATA <= x"f580";
            when "00" & x"a34" => DATA <= x"2001";
            when "00" & x"a35" => DATA <= x"e098";
            when "00" & x"a36" => DATA <= x"6100";
            when "00" & x"a37" => DATA <= x"f578";
            when "00" & x"a38" => DATA <= x"e198";
            when "00" & x"a39" => DATA <= x"6100";
            when "00" & x"a3a" => DATA <= x"f572";
            when "00" & x"a3b" => DATA <= x"7000";
            when "00" & x"a3c" => DATA <= x"6100";
            when "00" & x"a3d" => DATA <= x"f56c";
            when "00" & x"a3e" => DATA <= x"6100";
            when "00" & x"a3f" => DATA <= x"f568";
            when "00" & x"a40" => DATA <= x"6100";
            when "00" & x"a41" => DATA <= x"f564";
            when "00" & x"a42" => DATA <= x"221f";
            when "00" & x"a43" => DATA <= x"201f";
            when "00" & x"a44" => DATA <= x"023c";
            when "00" & x"a45" => DATA <= x"00fe";
            when "00" & x"a46" => DATA <= x"4e75";
            when "00" & x"a47" => DATA <= x"203c";
            when "00" & x"a48" => DATA <= x"003f";
            when "00" & x"a49" => DATA <= x"2d64";
            when "00" & x"a4a" => DATA <= x"003c";
            when "00" & x"a4b" => DATA <= x"0002";
            when "00" & x"a4c" => DATA <= x"4e75";
            when "00" & x"a4d" => DATA <= x"6100";
            when "00" & x"a4e" => DATA <= x"f584";
            when "00" & x"a4f" => DATA <= x"0000";
            when "00" & x"a50" => DATA <= x"0020";
            when "00" & x"a51" => DATA <= x"b03c";
            when "00" & x"a52" => DATA <= x"0079";
            when "00" & x"a53" => DATA <= x"4e75";
            when "00" & x"a54" => DATA <= x"2f0e";
            when "00" & x"a55" => DATA <= x"2f04";
            when "00" & x"a56" => DATA <= x"2c41";
            when "00" & x"a57" => DATA <= x"8643";
            when "00" & x"a58" => DATA <= x"6700";
            when "00" & x"a59" => DATA <= x"001e";
            when "00" & x"a5a" => DATA <= x"1816";
            when "00" & x"a5b" => DATA <= x"e144";
            when "00" & x"a5c" => DATA <= x"b940";
            when "00" & x"a5d" => DATA <= x"7807";
            when "00" & x"a5e" => DATA <= x"e340";
            when "00" & x"a5f" => DATA <= x"6400";
            when "00" & x"a60" => DATA <= x"0006";
            when "00" & x"a61" => DATA <= x"0a40";
            when "00" & x"a62" => DATA <= x"1021";
            when "00" & x"a63" => DATA <= x"51cc";
            when "00" & x"a64" => DATA <= x"fff4";
            when "00" & x"a65" => DATA <= x"dcc3";
            when "00" & x"a66" => DATA <= x"b48e";
            when "00" & x"a67" => DATA <= x"65e4";
            when "00" & x"a68" => DATA <= x"281f";
            when "00" & x"a69" => DATA <= x"2c5f";
            when "00" & x"a6a" => DATA <= x"023c";
            when "00" & x"a6b" => DATA <= x"00fd";
            when "00" & x"a6c" => DATA <= x"4e75";
            when "00" & x"a6d" => DATA <= x"1400";
            when "00" & x"a6e" => DATA <= x"708a";
            when "00" & x"a6f" => DATA <= x"7203";
            when "00" & x"a70" => DATA <= x"6100";
            when "00" & x"a71" => DATA <= x"f5f0";
            when "00" & x"a72" => DATA <= x"4e75";
            when "00" & x"a73" => DATA <= x"027c";
            when "00" & x"a74" => DATA <= x"dfff";
            when "00" & x"a75" => DATA <= x"4e75";
            when "00" & x"a76" => DATA <= x"b2bc";
            when "00" & x"a77" => DATA <= x"0000";
            when "00" & x"a78" => DATA <= x"00ff";
            when "00" & x"a79" => DATA <= x"6200";
            when "00" & x"a7a" => DATA <= x"0060";
            when "00" & x"a7b" => DATA <= x"2f08";
            when "00" & x"a7c" => DATA <= x"2040";
            when "00" & x"a7d" => DATA <= x"103c";
            when "00" & x"a7e" => DATA <= x"000a";
            when "00" & x"a7f" => DATA <= x"6100";
            when "00" & x"a80" => DATA <= x"eee2";
            when "00" & x"a81" => DATA <= x"1003";
            when "00" & x"a82" => DATA <= x"6100";
            when "00" & x"a83" => DATA <= x"eedc";
            when "00" & x"a84" => DATA <= x"1002";
            when "00" & x"a85" => DATA <= x"6100";
            when "00" & x"a86" => DATA <= x"eed6";
            when "00" & x"a87" => DATA <= x"1001";
            when "00" & x"a88" => DATA <= x"6100";
            when "00" & x"a89" => DATA <= x"eed0";
            when "00" & x"a8a" => DATA <= x"103c";
            when "00" & x"a8b" => DATA <= x"0007";
            when "00" & x"a8c" => DATA <= x"6100";
            when "00" & x"a8d" => DATA <= x"eec8";
            when "00" & x"a8e" => DATA <= x"103c";
            when "00" & x"a8f" => DATA <= x"0000";
            when "00" & x"a90" => DATA <= x"6100";
            when "00" & x"a91" => DATA <= x"eec0";
            when "00" & x"a92" => DATA <= x"6100";
            when "00" & x"a93" => DATA <= x"eeaa";
            when "00" & x"a94" => DATA <= x"b03c";
            when "00" & x"a95" => DATA <= x"0080";
            when "00" & x"a96" => DATA <= x"6700";
            when "00" & x"a97" => DATA <= x"001c";
            when "00" & x"a98" => DATA <= x"7200";
            when "00" & x"a99" => DATA <= x"6100";
            when "00" & x"a9a" => DATA <= x"ee9c";
            when "00" & x"a9b" => DATA <= x"10c0";
            when "00" & x"a9c" => DATA <= x"5241";
            when "00" & x"a9d" => DATA <= x"b03c";
            when "00" & x"a9e" => DATA <= x"000d";
            when "00" & x"a9f" => DATA <= x"66f2";
            when "00" & x"aa0" => DATA <= x"5341";
            when "00" & x"aa1" => DATA <= x"205f";
            when "00" & x"aa2" => DATA <= x"023c";
            when "00" & x"aa3" => DATA <= x"00fe";
            when "00" & x"aa4" => DATA <= x"4e75";
            when "00" & x"aa5" => DATA <= x"205f";
            when "00" & x"aa6" => DATA <= x"5341";
            when "00" & x"aa7" => DATA <= x"003c";
            when "00" & x"aa8" => DATA <= x"0001";
            when "00" & x"aa9" => DATA <= x"4e75";
            when "00" & x"aaa" => DATA <= x"003c";
            when "00" & x"aab" => DATA <= x"0002";
            when "00" & x"aac" => DATA <= x"4e75";
            when "00" & x"aad" => DATA <= x"2f03";
            when "00" & x"aae" => DATA <= x"2639";
            when "00" & x"aaf" => DATA <= x"003f";
            when "00" & x"ab0" => DATA <= x"3eda";
            when "00" & x"ab1" => DATA <= x"6100";
            when "00" & x"ab2" => DATA <= x"0006";
            when "00" & x"ab3" => DATA <= x"261f";
            when "00" & x"ab4" => DATA <= x"4e75";
            when "00" & x"ab5" => DATA <= x"2f0e";
            when "00" & x"ab6" => DATA <= x"2f0d";
            when "00" & x"ab7" => DATA <= x"2c41";
            when "00" & x"ab8" => DATA <= x"2a43";
            when "00" & x"ab9" => DATA <= x"101e";
            when "00" & x"aba" => DATA <= x"b03c";
            when "00" & x"abb" => DATA <= x"0025";
            when "00" & x"abc" => DATA <= x"6700";
            when "00" & x"abd" => DATA <= x"0010";
            when "00" & x"abe" => DATA <= x"1ac0";
            when "00" & x"abf" => DATA <= x"b03c";
            when "00" & x"ac0" => DATA <= x"0000";
            when "00" & x"ac1" => DATA <= x"66ee";
            when "00" & x"ac2" => DATA <= x"2a5f";
            when "00" & x"ac3" => DATA <= x"2c5f";
            when "00" & x"ac4" => DATA <= x"4e75";
            when "00" & x"ac5" => DATA <= x"101e";
            when "00" & x"ac6" => DATA <= x"b03c";
            when "00" & x"ac7" => DATA <= x"0030";
            when "00" & x"ac8" => DATA <= x"6600";
            when "00" & x"ac9" => DATA <= x"0008";
            when "00" & x"aca" => DATA <= x"1afc";
            when "00" & x"acb" => DATA <= x"0000";
            when "00" & x"acc" => DATA <= x"60d8";
            when "00" & x"acd" => DATA <= x"c03c";
            when "00" & x"ace" => DATA <= x"00df";
            when "00" & x"acf" => DATA <= x"b03c";
            when "00" & x"ad0" => DATA <= x"0025";
            when "00" & x"ad1" => DATA <= x"6600";
            when "00" & x"ad2" => DATA <= x"0008";
            when "00" & x"ad3" => DATA <= x"1afc";
            when "00" & x"ad4" => DATA <= x"0025";
            when "00" & x"ad5" => DATA <= x"60c6";
            when "00" & x"ad6" => DATA <= x"b03c";
            when "00" & x"ad7" => DATA <= x"005a";
            when "00" & x"ad8" => DATA <= x"6600";
            when "00" & x"ad9" => DATA <= x"0006";
            when "00" & x"ada" => DATA <= x"123c";
            when "00" & x"adb" => DATA <= x"005a";
            when "00" & x"adc" => DATA <= x"e158";
            when "00" & x"add" => DATA <= x"101e";
            when "00" & x"ade" => DATA <= x"c07c";
            when "00" & x"adf" => DATA <= x"dfdf";
            when "00" & x"ae0" => DATA <= x"b07c";
            when "00" & x"ae1" => DATA <= x"4353";
            when "00" & x"ae2" => DATA <= x"6700";
            when "00" & x"ae3" => DATA <= x"00aa";
            when "00" & x"ae4" => DATA <= x"b07c";
            when "00" & x"ae5" => DATA <= x"5345";
            when "00" & x"ae6" => DATA <= x"6700";
            when "00" & x"ae7" => DATA <= x"00a2";
            when "00" & x"ae8" => DATA <= x"b07c";
            when "00" & x"ae9" => DATA <= x"4d49";
            when "00" & x"aea" => DATA <= x"6700";
            when "00" & x"aeb" => DATA <= x"009a";
            when "00" & x"aec" => DATA <= x"b07c";
            when "00" & x"aed" => DATA <= x"3132";
            when "00" & x"aee" => DATA <= x"6700";
            when "00" & x"aef" => DATA <= x"0092";
            when "00" & x"af0" => DATA <= x"b07c";
            when "00" & x"af1" => DATA <= x"3234";
            when "00" & x"af2" => DATA <= x"6700";
            when "00" & x"af3" => DATA <= x"008a";
            when "00" & x"af4" => DATA <= x"b07c";
            when "00" & x"af5" => DATA <= x"414d";
            when "00" & x"af6" => DATA <= x"6700";
            when "00" & x"af7" => DATA <= x"0082";
            when "00" & x"af8" => DATA <= x"b07c";
            when "00" & x"af9" => DATA <= x"504d";
            when "00" & x"afa" => DATA <= x"6700";
            when "00" & x"afb" => DATA <= x"007a";
            when "00" & x"afc" => DATA <= x"b07c";
            when "00" & x"afd" => DATA <= x"5745";
            when "00" & x"afe" => DATA <= x"6700";
            when "00" & x"aff" => DATA <= x"0072";
            when "00" & x"b00" => DATA <= x"b07c";
            when "00" & x"b01" => DATA <= x"5733";
            when "00" & x"b02" => DATA <= x"6700";
            when "00" & x"b03" => DATA <= x"006a";
            when "00" & x"b04" => DATA <= x"b07c";
            when "00" & x"b05" => DATA <= x"574e";
            when "00" & x"b06" => DATA <= x"6700";
            when "00" & x"b07" => DATA <= x"0062";
            when "00" & x"b08" => DATA <= x"b07c";
            when "00" & x"b09" => DATA <= x"4459";
            when "00" & x"b0a" => DATA <= x"6700";
            when "00" & x"b0b" => DATA <= x"005a";
            when "00" & x"b0c" => DATA <= x"b07c";
            when "00" & x"b0d" => DATA <= x"5354";
            when "00" & x"b0e" => DATA <= x"6700";
            when "00" & x"b0f" => DATA <= x"0052";
            when "00" & x"b10" => DATA <= x"b07c";
            when "00" & x"b11" => DATA <= x"4d4f";
            when "00" & x"b12" => DATA <= x"6700";
            when "00" & x"b13" => DATA <= x"004a";
            when "00" & x"b14" => DATA <= x"b07c";
            when "00" & x"b15" => DATA <= x"4d33";
            when "00" & x"b16" => DATA <= x"6700";
            when "00" & x"b17" => DATA <= x"0042";
            when "00" & x"b18" => DATA <= x"b07c";
            when "00" & x"b19" => DATA <= x"4d4e";
            when "00" & x"b1a" => DATA <= x"6700";
            when "00" & x"b1b" => DATA <= x"003a";
            when "00" & x"b1c" => DATA <= x"b07c";
            when "00" & x"b1d" => DATA <= x"4345";
            when "00" & x"b1e" => DATA <= x"6700";
            when "00" & x"b1f" => DATA <= x"0032";
            when "00" & x"b20" => DATA <= x"b07c";
            when "00" & x"b21" => DATA <= x"5952";
            when "00" & x"b22" => DATA <= x"6700";
            when "00" & x"b23" => DATA <= x"002a";
            when "00" & x"b24" => DATA <= x"b07c";
            when "00" & x"b25" => DATA <= x"574b";
            when "00" & x"b26" => DATA <= x"6700";
            when "00" & x"b27" => DATA <= x"0022";
            when "00" & x"b28" => DATA <= x"b07c";
            when "00" & x"b29" => DATA <= x"444e";
            when "00" & x"b2a" => DATA <= x"6700";
            when "00" & x"b2b" => DATA <= x"001a";
            when "00" & x"b2c" => DATA <= x"b07c";
            when "00" & x"b2d" => DATA <= x"545a";
            when "00" & x"b2e" => DATA <= x"6700";
            when "00" & x"b2f" => DATA <= x"0012";
            when "00" & x"b30" => DATA <= x"2a5f";
            when "00" & x"b31" => DATA <= x"2c5f";
            when "00" & x"b32" => DATA <= x"203c";
            when "00" & x"b33" => DATA <= x"003f";
            when "00" & x"b34" => DATA <= x"2eac";
            when "00" & x"b35" => DATA <= x"003c";
            when "00" & x"b36" => DATA <= x"0002";
            when "00" & x"b37" => DATA <= x"4e75";
            when "00" & x"b38" => DATA <= x"6000";
            when "00" & x"b39" => DATA <= x"ff00";
            when "00" & x"b3a" => DATA <= x"b4bc";
            when "00" & x"b3b" => DATA <= x"0000";
            when "00" & x"b3c" => DATA <= x"0002";
            when "00" & x"b3d" => DATA <= x"6f00";
            when "00" & x"b3e" => DATA <= x"0484";
            when "00" & x"b3f" => DATA <= x"5582";
            when "00" & x"b40" => DATA <= x"2f0e";
            when "00" & x"b41" => DATA <= x"48e7";
            when "00" & x"b42" => DATA <= x"7000";
            when "00" & x"b43" => DATA <= x"343c";
            when "00" & x"b44" => DATA <= x"0000";
            when "00" & x"b45" => DATA <= x"e898";
            when "00" & x"b46" => DATA <= x"6000";
            when "00" & x"b47" => DATA <= x"0072";
            when "00" & x"b48" => DATA <= x"b4bc";
            when "00" & x"b49" => DATA <= x"0000";
            when "00" & x"b4a" => DATA <= x"0003";
            when "00" & x"b4b" => DATA <= x"6f00";
            when "00" & x"b4c" => DATA <= x"0468";
            when "00" & x"b4d" => DATA <= x"5782";
            when "00" & x"b4e" => DATA <= x"2f0e";
            when "00" & x"b4f" => DATA <= x"48e7";
            when "00" & x"b50" => DATA <= x"7000";
            when "00" & x"b51" => DATA <= x"343c";
            when "00" & x"b52" => DATA <= x"0001";
            when "00" & x"b53" => DATA <= x"e098";
            when "00" & x"b54" => DATA <= x"6000";
            when "00" & x"b55" => DATA <= x"0056";
            when "00" & x"b56" => DATA <= x"b4bc";
            when "00" & x"b57" => DATA <= x"0000";
            when "00" & x"b58" => DATA <= x"0005";
            when "00" & x"b59" => DATA <= x"6f00";
            when "00" & x"b5a" => DATA <= x"044c";
            when "00" & x"b5b" => DATA <= x"5b82";
            when "00" & x"b5c" => DATA <= x"2f0e";
            when "00" & x"b5d" => DATA <= x"48e7";
            when "00" & x"b5e" => DATA <= x"7000";
            when "00" & x"b5f" => DATA <= x"343c";
            when "00" & x"b60" => DATA <= x"0003";
            when "00" & x"b61" => DATA <= x"e198";
            when "00" & x"b62" => DATA <= x"e198";
            when "00" & x"b63" => DATA <= x"6000";
            when "00" & x"b64" => DATA <= x"0038";
            when "00" & x"b65" => DATA <= x"b4bc";
            when "00" & x"b66" => DATA <= x"0000";
            when "00" & x"b67" => DATA <= x"0007";
            when "00" & x"b68" => DATA <= x"6f00";
            when "00" & x"b69" => DATA <= x"042e";
            when "00" & x"b6a" => DATA <= x"5f82";
            when "00" & x"b6b" => DATA <= x"2f0e";
            when "00" & x"b6c" => DATA <= x"48e7";
            when "00" & x"b6d" => DATA <= x"7000";
            when "00" & x"b6e" => DATA <= x"343c";
            when "00" & x"b6f" => DATA <= x"0005";
            when "00" & x"b70" => DATA <= x"e098";
            when "00" & x"b71" => DATA <= x"6000";
            when "00" & x"b72" => DATA <= x"001c";
            when "00" & x"b73" => DATA <= x"b4bc";
            when "00" & x"b74" => DATA <= x"0000";
            when "00" & x"b75" => DATA <= x"0009";
            when "00" & x"b76" => DATA <= x"6f00";
            when "00" & x"b77" => DATA <= x"0412";
            when "00" & x"b78" => DATA <= x"0482";
            when "00" & x"b79" => DATA <= x"0000";
            when "00" & x"b7a" => DATA <= x"0009";
            when "00" & x"b7b" => DATA <= x"2f0e";
            when "00" & x"b7c" => DATA <= x"48e7";
            when "00" & x"b7d" => DATA <= x"7000";
            when "00" & x"b7e" => DATA <= x"343c";
            when "00" & x"b7f" => DATA <= x"0007";
            when "00" & x"b80" => DATA <= x"2c41";
            when "00" & x"b81" => DATA <= x"2200";
            when "00" & x"b82" => DATA <= x"e999";
            when "00" & x"b83" => DATA <= x"1001";
            when "00" & x"b84" => DATA <= x"c03c";
            when "00" & x"b85" => DATA <= x"000f";
            when "00" & x"b86" => DATA <= x"163c";
            when "00" & x"b87" => DATA <= x"0009";
            when "00" & x"b88" => DATA <= x"9600";
            when "00" & x"b89" => DATA <= x"0600";
            when "00" & x"b8a" => DATA <= x"0030";
            when "00" & x"b8b" => DATA <= x"0c00";
            when "00" & x"b8c" => DATA <= x"003a";
            when "00" & x"b8d" => DATA <= x"6500";
            when "00" & x"b8e" => DATA <= x"0004";
            when "00" & x"b8f" => DATA <= x"5e00";
            when "00" & x"b90" => DATA <= x"1cc0";
            when "00" & x"b91" => DATA <= x"51ca";
            when "00" & x"b92" => DATA <= x"ffe0";
            when "00" & x"b93" => DATA <= x"1cbc";
            when "00" & x"b94" => DATA <= x"0000";
            when "00" & x"b95" => DATA <= x"4cdf";
            when "00" & x"b96" => DATA <= x"000e";
            when "00" & x"b97" => DATA <= x"2001";
            when "00" & x"b98" => DATA <= x"220e";
            when "00" & x"b99" => DATA <= x"2c5f";
            when "00" & x"b9a" => DATA <= x"023c";
            when "00" & x"b9b" => DATA <= x"00fd";
            when "00" & x"b9c" => DATA <= x"4e75";
            when "00" & x"b9d" => DATA <= x"003c";
            when "00" & x"b9e" => DATA <= x"0002";
            when "00" & x"b9f" => DATA <= x"4e75";
            when "00" & x"ba0" => DATA <= x"b4bc";
            when "00" & x"ba1" => DATA <= x"0000";
            when "00" & x"ba2" => DATA <= x"0004";
            when "00" & x"ba3" => DATA <= x"6500";
            when "00" & x"ba4" => DATA <= x"03b8";
            when "00" & x"ba5" => DATA <= x"b0bc";
            when "00" & x"ba6" => DATA <= x"0000";
            when "00" & x"ba7" => DATA <= x"0100";
            when "00" & x"ba8" => DATA <= x"6400";
            when "00" & x"ba9" => DATA <= x"01b2";
            when "00" & x"baa" => DATA <= x"7c03";
            when "00" & x"bab" => DATA <= x"6000";
            when "00" & x"bac" => DATA <= x"0042";
            when "00" & x"bad" => DATA <= x"b4bc";
            when "00" & x"bae" => DATA <= x"0000";
            when "00" & x"baf" => DATA <= x"0006";
            when "00" & x"bb0" => DATA <= x"6500";
            when "00" & x"bb1" => DATA <= x"039e";
            when "00" & x"bb2" => DATA <= x"b0bc";
            when "00" & x"bb3" => DATA <= x"0001";
            when "00" & x"bb4" => DATA <= x"0000";
            when "00" & x"bb5" => DATA <= x"6400";
            when "00" & x"bb6" => DATA <= x"0198";
            when "00" & x"bb7" => DATA <= x"7c05";
            when "00" & x"bb8" => DATA <= x"6000";
            when "00" & x"bb9" => DATA <= x"0028";
            when "00" & x"bba" => DATA <= x"b4bc";
            when "00" & x"bbb" => DATA <= x"0000";
            when "00" & x"bbc" => DATA <= x"0009";
            when "00" & x"bbd" => DATA <= x"6500";
            when "00" & x"bbe" => DATA <= x"0384";
            when "00" & x"bbf" => DATA <= x"b0bc";
            when "00" & x"bc0" => DATA <= x"0100";
            when "00" & x"bc1" => DATA <= x"0000";
            when "00" & x"bc2" => DATA <= x"6400";
            when "00" & x"bc3" => DATA <= x"017e";
            when "00" & x"bc4" => DATA <= x"7c08";
            when "00" & x"bc5" => DATA <= x"6000";
            when "00" & x"bc6" => DATA <= x"000e";
            when "00" & x"bc7" => DATA <= x"b4bc";
            when "00" & x"bc8" => DATA <= x"0000";
            when "00" & x"bc9" => DATA <= x"000b";
            when "00" & x"bca" => DATA <= x"6500";
            when "00" & x"bcb" => DATA <= x"036a";
            when "00" & x"bcc" => DATA <= x"7c0a";
            when "00" & x"bcd" => DATA <= x"c38d";
            when "00" & x"bce" => DATA <= x"48e7";
            when "00" & x"bcf" => DATA <= x"ff00";
            when "00" & x"bd0" => DATA <= x"2e00";
            when "00" & x"bd1" => DATA <= x"6700";
            when "00" & x"bd2" => DATA <= x"0058";
            when "00" & x"bd3" => DATA <= x"6000";
            when "00" & x"bd4" => DATA <= x"0002";
            when "00" & x"bd5" => DATA <= x"4244";
            when "00" & x"bd6" => DATA <= x"7401";
            when "00" & x"bd7" => DATA <= x"2206";
            when "00" & x"bd8" => DATA <= x"5381";
            when "00" & x"bd9" => DATA <= x"6700";
            when "00" & x"bda" => DATA <= x"001c";
            when "00" & x"bdb" => DATA <= x"3602";
            when "00" & x"bdc" => DATA <= x"c6fc";
            when "00" & x"bdd" => DATA <= x"000a";
            when "00" & x"bde" => DATA <= x"4842";
            when "00" & x"bdf" => DATA <= x"c4fc";
            when "00" & x"be0" => DATA <= x"000a";
            when "00" & x"be1" => DATA <= x"4843";
            when "00" & x"be2" => DATA <= x"d443";
            when "00" & x"be3" => DATA <= x"4842";
            when "00" & x"be4" => DATA <= x"4843";
            when "00" & x"be5" => DATA <= x"3403";
            when "00" & x"be6" => DATA <= x"5381";
            when "00" & x"be7" => DATA <= x"66e6";
            when "00" & x"be8" => DATA <= x"4280";
            when "00" & x"be9" => DATA <= x"be82";
            when "00" & x"bea" => DATA <= x"6500";
            when "00" & x"beb" => DATA <= x"0008";
            when "00" & x"bec" => DATA <= x"5280";
            when "00" & x"bed" => DATA <= x"9e82";
            when "00" & x"bee" => DATA <= x"60f4";
            when "00" & x"bef" => DATA <= x"4a00";
            when "00" & x"bf0" => DATA <= x"6600";
            when "00" & x"bf1" => DATA <= x"0008";
            when "00" & x"bf2" => DATA <= x"4a44";
            when "00" & x"bf3" => DATA <= x"6700";
            when "00" & x"bf4" => DATA <= x"000a";
            when "00" & x"bf5" => DATA <= x"0600";
            when "00" & x"bf6" => DATA <= x"0030";
            when "00" & x"bf7" => DATA <= x"1ac0";
            when "00" & x"bf8" => DATA <= x"1800";
            when "00" & x"bf9" => DATA <= x"5386";
            when "00" & x"bfa" => DATA <= x"66b6";
            when "00" & x"bfb" => DATA <= x"4a44";
            when "00" & x"bfc" => DATA <= x"6600";
            when "00" & x"bfd" => DATA <= x"0006";
            when "00" & x"bfe" => DATA <= x"1afc";
            when "00" & x"bff" => DATA <= x"0030";
            when "00" & x"c00" => DATA <= x"1abc";
            when "00" & x"c01" => DATA <= x"0000";
            when "00" & x"c02" => DATA <= x"4cdf";
            when "00" & x"c03" => DATA <= x"00ff";
            when "00" & x"c04" => DATA <= x"c38d";
            when "00" & x"c05" => DATA <= x"023c";
            when "00" & x"c06" => DATA <= x"00fd";
            when "00" & x"c07" => DATA <= x"4e75";
            when "00" & x"c08" => DATA <= x"b4bc";
            when "00" & x"c09" => DATA <= x"0000";
            when "00" & x"c0a" => DATA <= x"0005";
            when "00" & x"c0b" => DATA <= x"6500";
            when "00" & x"c0c" => DATA <= x"02e8";
            when "00" & x"c0d" => DATA <= x"b0bc";
            when "00" & x"c0e" => DATA <= x"0000";
            when "00" & x"c0f" => DATA <= x"0100";
            when "00" & x"c10" => DATA <= x"6400";
            when "00" & x"c11" => DATA <= x"00e2";
            when "00" & x"c12" => DATA <= x"0800";
            when "00" & x"c13" => DATA <= x"0007";
            when "00" & x"c14" => DATA <= x"6700";
            when "00" & x"c15" => DATA <= x"0008";
            when "00" & x"c16" => DATA <= x"0080";
            when "00" & x"c17" => DATA <= x"ffff";
            when "00" & x"c18" => DATA <= x"ff00";
            when "00" & x"c19" => DATA <= x"7c03";
            when "00" & x"c1a" => DATA <= x"6000";
            when "00" & x"c1b" => DATA <= x"005e";
            when "00" & x"c1c" => DATA <= x"b4bc";
            when "00" & x"c1d" => DATA <= x"0000";
            when "00" & x"c1e" => DATA <= x"0007";
            when "00" & x"c1f" => DATA <= x"6500";
            when "00" & x"c20" => DATA <= x"02c0";
            when "00" & x"c21" => DATA <= x"b0bc";
            when "00" & x"c22" => DATA <= x"0001";
            when "00" & x"c23" => DATA <= x"0000";
            when "00" & x"c24" => DATA <= x"6400";
            when "00" & x"c25" => DATA <= x"00ba";
            when "00" & x"c26" => DATA <= x"0800";
            when "00" & x"c27" => DATA <= x"000f";
            when "00" & x"c28" => DATA <= x"6700";
            when "00" & x"c29" => DATA <= x"0008";
            when "00" & x"c2a" => DATA <= x"0080";
            when "00" & x"c2b" => DATA <= x"ffff";
            when "00" & x"c2c" => DATA <= x"0000";
            when "00" & x"c2d" => DATA <= x"7c05";
            when "00" & x"c2e" => DATA <= x"6000";
            when "00" & x"c2f" => DATA <= x"0036";
            when "00" & x"c30" => DATA <= x"b4bc";
            when "00" & x"c31" => DATA <= x"0000";
            when "00" & x"c32" => DATA <= x"000b";
            when "00" & x"c33" => DATA <= x"6500";
            when "00" & x"c34" => DATA <= x"0298";
            when "00" & x"c35" => DATA <= x"b0bc";
            when "00" & x"c36" => DATA <= x"0100";
            when "00" & x"c37" => DATA <= x"0000";
            when "00" & x"c38" => DATA <= x"6400";
            when "00" & x"c39" => DATA <= x"0092";
            when "00" & x"c3a" => DATA <= x"0800";
            when "00" & x"c3b" => DATA <= x"0017";
            when "00" & x"c3c" => DATA <= x"6700";
            when "00" & x"c3d" => DATA <= x"0008";
            when "00" & x"c3e" => DATA <= x"0080";
            when "00" & x"c3f" => DATA <= x"ff00";
            when "00" & x"c40" => DATA <= x"0000";
            when "00" & x"c41" => DATA <= x"7c08";
            when "00" & x"c42" => DATA <= x"6000";
            when "00" & x"c43" => DATA <= x"000e";
            when "00" & x"c44" => DATA <= x"b4bc";
            when "00" & x"c45" => DATA <= x"0000";
            when "00" & x"c46" => DATA <= x"000d";
            when "00" & x"c47" => DATA <= x"6500";
            when "00" & x"c48" => DATA <= x"0270";
            when "00" & x"c49" => DATA <= x"7c0a";
            when "00" & x"c4a" => DATA <= x"c38d";
            when "00" & x"c4b" => DATA <= x"48e7";
            when "00" & x"c4c" => DATA <= x"ff00";
            when "00" & x"c4d" => DATA <= x"2e00";
            when "00" & x"c4e" => DATA <= x"6a08";
            when "00" & x"c4f" => DATA <= x"4487";
            when "00" & x"c50" => DATA <= x"6b4e";
            when "00" & x"c51" => DATA <= x"1afc";
            when "00" & x"c52" => DATA <= x"002d";
            when "00" & x"c53" => DATA <= x"4244";
            when "00" & x"c54" => DATA <= x"7a01";
            when "00" & x"c55" => DATA <= x"2206";
            when "00" & x"c56" => DATA <= x"5381";
            when "00" & x"c57" => DATA <= x"671a";
            when "00" & x"c58" => DATA <= x"3605";
            when "00" & x"c59" => DATA <= x"c6fc";
            when "00" & x"c5a" => DATA <= x"000a";
            when "00" & x"c5b" => DATA <= x"4845";
            when "00" & x"c5c" => DATA <= x"cafc";
            when "00" & x"c5d" => DATA <= x"000a";
            when "00" & x"c5e" => DATA <= x"4843";
            when "00" & x"c5f" => DATA <= x"da43";
            when "00" & x"c60" => DATA <= x"4845";
            when "00" & x"c61" => DATA <= x"4843";
            when "00" & x"c62" => DATA <= x"3a03";
            when "00" & x"c63" => DATA <= x"5381";
            when "00" & x"c64" => DATA <= x"66e6";
            when "00" & x"c65" => DATA <= x"4280";
            when "00" & x"c66" => DATA <= x"be85";
            when "00" & x"c67" => DATA <= x"6d06";
            when "00" & x"c68" => DATA <= x"5280";
            when "00" & x"c69" => DATA <= x"9e85";
            when "00" & x"c6a" => DATA <= x"60f6";
            when "00" & x"c6b" => DATA <= x"4a00";
            when "00" & x"c6c" => DATA <= x"6604";
            when "00" & x"c6d" => DATA <= x"4a44";
            when "00" & x"c6e" => DATA <= x"6708";
            when "00" & x"c6f" => DATA <= x"0600";
            when "00" & x"c70" => DATA <= x"0030";
            when "00" & x"c71" => DATA <= x"1ac0";
            when "00" & x"c72" => DATA <= x"1800";
            when "00" & x"c73" => DATA <= x"5386";
            when "00" & x"c74" => DATA <= x"66be";
            when "00" & x"c75" => DATA <= x"4a44";
            when "00" & x"c76" => DATA <= x"6600";
            when "00" & x"c77" => DATA <= x"0006";
            when "00" & x"c78" => DATA <= x"1afc";
            when "00" & x"c79" => DATA <= x"0030";
            when "00" & x"c7a" => DATA <= x"1abc";
            when "00" & x"c7b" => DATA <= x"0000";
            when "00" & x"c7c" => DATA <= x"4cdf";
            when "00" & x"c7d" => DATA <= x"00ff";
            when "00" & x"c7e" => DATA <= x"c38d";
            when "00" & x"c7f" => DATA <= x"023c";
            when "00" & x"c80" => DATA <= x"00fd";
            when "00" & x"c81" => DATA <= x"4e75";
            when "00" & x"c82" => DATA <= x"003c";
            when "00" & x"c83" => DATA <= x"0002";
            when "00" & x"c84" => DATA <= x"4e75";
            when "00" & x"c85" => DATA <= x"b4bc";
            when "00" & x"c86" => DATA <= x"0000";
            when "00" & x"c87" => DATA <= x"0009";
            when "00" & x"c88" => DATA <= x"6f00";
            when "00" & x"c89" => DATA <= x"01ee";
            when "00" & x"c8a" => DATA <= x"0482";
            when "00" & x"c8b" => DATA <= x"0000";
            when "00" & x"c8c" => DATA <= x"0009";
            when "00" & x"c8d" => DATA <= x"2f0e";
            when "00" & x"c8e" => DATA <= x"48e7";
            when "00" & x"c8f" => DATA <= x"7000";
            when "00" & x"c90" => DATA <= x"7407";
            when "00" & x"c91" => DATA <= x"e098";
            when "00" & x"c92" => DATA <= x"6000";
            when "00" & x"c93" => DATA <= x"0058";
            when "00" & x"c94" => DATA <= x"b4bc";
            when "00" & x"c95" => DATA <= x"0000";
            when "00" & x"c96" => DATA <= x"0011";
            when "00" & x"c97" => DATA <= x"6f00";
            when "00" & x"c98" => DATA <= x"01d0";
            when "00" & x"c99" => DATA <= x"0482";
            when "00" & x"c9a" => DATA <= x"0000";
            when "00" & x"c9b" => DATA <= x"0011";
            when "00" & x"c9c" => DATA <= x"2f0e";
            when "00" & x"c9d" => DATA <= x"48e7";
            when "00" & x"c9e" => DATA <= x"7000";
            when "00" & x"c9f" => DATA <= x"740f";
            when "00" & x"ca0" => DATA <= x"e198";
            when "00" & x"ca1" => DATA <= x"e198";
            when "00" & x"ca2" => DATA <= x"6000";
            when "00" & x"ca3" => DATA <= x"0038";
            when "00" & x"ca4" => DATA <= x"b4bc";
            when "00" & x"ca5" => DATA <= x"0000";
            when "00" & x"ca6" => DATA <= x"0019";
            when "00" & x"ca7" => DATA <= x"6f00";
            when "00" & x"ca8" => DATA <= x"01b0";
            when "00" & x"ca9" => DATA <= x"0482";
            when "00" & x"caa" => DATA <= x"0000";
            when "00" & x"cab" => DATA <= x"0019";
            when "00" & x"cac" => DATA <= x"2f0e";
            when "00" & x"cad" => DATA <= x"48e7";
            when "00" & x"cae" => DATA <= x"7000";
            when "00" & x"caf" => DATA <= x"7417";
            when "00" & x"cb0" => DATA <= x"e098";
            when "00" & x"cb1" => DATA <= x"6000";
            when "00" & x"cb2" => DATA <= x"001a";
            when "00" & x"cb3" => DATA <= x"b4bc";
            when "00" & x"cb4" => DATA <= x"0000";
            when "00" & x"cb5" => DATA <= x"0021";
            when "00" & x"cb6" => DATA <= x"6f00";
            when "00" & x"cb7" => DATA <= x"0192";
            when "00" & x"cb8" => DATA <= x"0482";
            when "00" & x"cb9" => DATA <= x"0000";
            when "00" & x"cba" => DATA <= x"0021";
            when "00" & x"cbb" => DATA <= x"2f0e";
            when "00" & x"cbc" => DATA <= x"48e7";
            when "00" & x"cbd" => DATA <= x"7000";
            when "00" & x"cbe" => DATA <= x"741f";
            when "00" & x"cbf" => DATA <= x"2c41";
            when "00" & x"cc0" => DATA <= x"7600";
            when "00" & x"cc1" => DATA <= x"7230";
            when "00" & x"cc2" => DATA <= x"e380";
            when "00" & x"cc3" => DATA <= x"c303";
            when "00" & x"cc4" => DATA <= x"1cc1";
            when "00" & x"cc5" => DATA <= x"51ca";
            when "00" & x"cc6" => DATA <= x"fff6";
            when "00" & x"cc7" => DATA <= x"1cbc";
            when "00" & x"cc8" => DATA <= x"0000";
            when "00" & x"cc9" => DATA <= x"4cdf";
            when "00" & x"cca" => DATA <= x"000e";
            when "00" & x"ccb" => DATA <= x"2001";
            when "00" & x"ccc" => DATA <= x"220e";
            when "00" & x"ccd" => DATA <= x"2c5f";
            when "00" & x"cce" => DATA <= x"023c";
            when "00" & x"ccf" => DATA <= x"00fd";
            when "00" & x"cd0" => DATA <= x"4e75";
            when "00" & x"cd1" => DATA <= x"6100";
            when "00" & x"cd2" => DATA <= x"fe6c";
            when "00" & x"cd3" => DATA <= x"2f07";
            when "00" & x"cd4" => DATA <= x"7e05";
            when "00" & x"cd5" => DATA <= x"6100";
            when "00" & x"cd6" => DATA <= x"0122";
            when "00" & x"cd7" => DATA <= x"2e1f";
            when "00" & x"cd8" => DATA <= x"4e75";
            when "00" & x"cd9" => DATA <= x"6100";
            when "00" & x"cda" => DATA <= x"fe84";
            when "00" & x"cdb" => DATA <= x"2f07";
            when "00" & x"cdc" => DATA <= x"7e07";
            when "00" & x"cdd" => DATA <= x"6100";
            when "00" & x"cde" => DATA <= x"0112";
            when "00" & x"cdf" => DATA <= x"2e1f";
            when "00" & x"ce0" => DATA <= x"4e75";
            when "00" & x"ce1" => DATA <= x"6100";
            when "00" & x"ce2" => DATA <= x"fe9c";
            when "00" & x"ce3" => DATA <= x"2f07";
            when "00" & x"ce4" => DATA <= x"7e09";
            when "00" & x"ce5" => DATA <= x"6100";
            when "00" & x"ce6" => DATA <= x"0102";
            when "00" & x"ce7" => DATA <= x"2e1f";
            when "00" & x"ce8" => DATA <= x"4e75";
            when "00" & x"ce9" => DATA <= x"6100";
            when "00" & x"cea" => DATA <= x"feb4";
            when "00" & x"ceb" => DATA <= x"2f07";
            when "00" & x"cec" => DATA <= x"7e0c";
            when "00" & x"ced" => DATA <= x"6100";
            when "00" & x"cee" => DATA <= x"00f2";
            when "00" & x"cef" => DATA <= x"2e1f";
            when "00" & x"cf0" => DATA <= x"4e75";
            when "00" & x"cf1" => DATA <= x"2f01";
            when "00" & x"cf2" => DATA <= x"2f06";
            when "00" & x"cf3" => DATA <= x"2f07";
            when "00" & x"cf4" => DATA <= x"2f0e";
            when "00" & x"cf5" => DATA <= x"2c40";
            when "00" & x"cf6" => DATA <= x"2c1e";
            when "00" & x"cf7" => DATA <= x"2e1e";
            when "00" & x"cf8" => DATA <= x"0c87";
            when "00" & x"cf9" => DATA <= x"0000";
            when "00" & x"cfa" => DATA <= x"0100";
            when "00" & x"cfb" => DATA <= x"6400";
            when "00" & x"cfc" => DATA <= x"003a";
            when "00" & x"cfd" => DATA <= x"0c86";
            when "00" & x"cfe" => DATA <= x"0000";
            when "00" & x"cff" => DATA <= x"0100";
            when "00" & x"d00" => DATA <= x"6400";
            when "00" & x"d01" => DATA <= x"003e";
            when "00" & x"d02" => DATA <= x"4a47";
            when "00" & x"d03" => DATA <= x"6700";
            when "00" & x"d04" => DATA <= x"0016";
            when "00" & x"d05" => DATA <= x"1007";
            when "00" & x"d06" => DATA <= x"6100";
            when "00" & x"d07" => DATA <= x"fd32";
            when "00" & x"d08" => DATA <= x"4a41";
            when "00" & x"d09" => DATA <= x"6700";
            when "00" & x"d0a" => DATA <= x"00ec";
            when "00" & x"d0b" => DATA <= x"2c41";
            when "00" & x"d0c" => DATA <= x"1cfc";
            when "00" & x"d0d" => DATA <= x"002e";
            when "00" & x"d0e" => DATA <= x"220e";
            when "00" & x"d0f" => DATA <= x"1006";
            when "00" & x"d10" => DATA <= x"6100";
            when "00" & x"d11" => DATA <= x"fd1e";
            when "00" & x"d12" => DATA <= x"2c5f";
            when "00" & x"d13" => DATA <= x"2e1f";
            when "00" & x"d14" => DATA <= x"2c1f";
            when "00" & x"d15" => DATA <= x"201f";
            when "00" & x"d16" => DATA <= x"023c";
            when "00" & x"d17" => DATA <= x"00fd";
            when "00" & x"d18" => DATA <= x"4e75";
            when "00" & x"d19" => DATA <= x"2f7c";
            when "00" & x"d1a" => DATA <= x"003f";
            when "00" & x"d1b" => DATA <= x"2edc";
            when "00" & x"d1c" => DATA <= x"000c";
            when "00" & x"d1d" => DATA <= x"003c";
            when "00" & x"d1e" => DATA <= x"0002";
            when "00" & x"d1f" => DATA <= x"60e4";
            when "00" & x"d20" => DATA <= x"2f7c";
            when "00" & x"d21" => DATA <= x"003f";
            when "00" & x"d22" => DATA <= x"2ec4";
            when "00" & x"d23" => DATA <= x"000c";
            when "00" & x"d24" => DATA <= x"003c";
            when "00" & x"d25" => DATA <= x"0002";
            when "00" & x"d26" => DATA <= x"60d6";
            when "00" & x"d27" => DATA <= x"2f07";
            when "00" & x"d28" => DATA <= x"2f01";
            when "00" & x"d29" => DATA <= x"2200";
            when "00" & x"d2a" => DATA <= x"0281";
            when "00" & x"d2b" => DATA <= x"c000";
            when "00" & x"d2c" => DATA <= x"0000";
            when "00" & x"d2d" => DATA <= x"6700";
            when "00" & x"d2e" => DATA <= x"0014";
            when "00" & x"d2f" => DATA <= x"e089";
            when "00" & x"d30" => DATA <= x"e089";
            when "00" & x"d31" => DATA <= x"e089";
            when "00" & x"d32" => DATA <= x"ec89";
            when "00" & x"d33" => DATA <= x"2001";
            when "00" & x"d34" => DATA <= x"1e38";
            when "00" & x"d35" => DATA <= x"004d";
            when "00" & x"d36" => DATA <= x"6000";
            when "00" & x"d37" => DATA <= x"0034";
            when "00" & x"d38" => DATA <= x"2200";
            when "00" & x"d39" => DATA <= x"0281";
            when "00" & x"d3a" => DATA <= x"fff0";
            when "00" & x"d3b" => DATA <= x"0000";
            when "00" & x"d3c" => DATA <= x"6700";
            when "00" & x"d3d" => DATA <= x"0012";
            when "00" & x"d3e" => DATA <= x"e089";
            when "00" & x"d3f" => DATA <= x"e089";
            when "00" & x"d40" => DATA <= x"e889";
            when "00" & x"d41" => DATA <= x"2001";
            when "00" & x"d42" => DATA <= x"1e38";
            when "00" & x"d43" => DATA <= x"004b";
            when "00" & x"d44" => DATA <= x"6000";
            when "00" & x"d45" => DATA <= x"0018";
            when "00" & x"d46" => DATA <= x"2200";
            when "00" & x"d47" => DATA <= x"0281";
            when "00" & x"d48" => DATA <= x"ffff";
            when "00" & x"d49" => DATA <= x"fc00";
            when "00" & x"d4a" => DATA <= x"6700";
            when "00" & x"d4b" => DATA <= x"000c";
            when "00" & x"d4c" => DATA <= x"e089";
            when "00" & x"d4d" => DATA <= x"e489";
            when "00" & x"d4e" => DATA <= x"2001";
            when "00" & x"d4f" => DATA <= x"1e3c";
            when "00" & x"d50" => DATA <= x"0000";
            when "00" & x"d51" => DATA <= x"221f";
            when "00" & x"d52" => DATA <= x"6100";
            when "00" & x"d53" => DATA <= x"fce8";
            when "00" & x"d54" => DATA <= x"2c41";
            when "00" & x"d55" => DATA <= x"1cfc";
            when "00" & x"d56" => DATA <= x"0020";
            when "00" & x"d57" => DATA <= x"1cc7";
            when "00" & x"d58" => DATA <= x"1cfc";
            when "00" & x"d59" => DATA <= x"0062";
            when "00" & x"d5a" => DATA <= x"1cfc";
            when "00" & x"d5b" => DATA <= x"0079";
            when "00" & x"d5c" => DATA <= x"1cfc";
            when "00" & x"d5d" => DATA <= x"0074";
            when "00" & x"d5e" => DATA <= x"1cfc";
            when "00" & x"d5f" => DATA <= x"0065";
            when "00" & x"d60" => DATA <= x"1cfc";
            when "00" & x"d61" => DATA <= x"0073";
            when "00" & x"d62" => DATA <= x"1cfc";
            when "00" & x"d63" => DATA <= x"0000";
            when "00" & x"d64" => DATA <= x"023c";
            when "00" & x"d65" => DATA <= x"00fd";
            when "00" & x"d66" => DATA <= x"4e75";
            when "00" & x"d67" => DATA <= x"2f0e";
            when "00" & x"d68" => DATA <= x"2f00";
            when "00" & x"d69" => DATA <= x"2f01";
            when "00" & x"d6a" => DATA <= x"2c40";
            when "00" & x"d6b" => DATA <= x"9280";
            when "00" & x"d6c" => DATA <= x"1dbc";
            when "00" & x"d6d" => DATA <= x"0000";
            when "00" & x"d6e" => DATA <= x"7000";
            when "00" & x"d6f" => DATA <= x"5387";
            when "00" & x"d70" => DATA <= x"1db6";
            when "00" & x"d71" => DATA <= x"1000";
            when "00" & x"d72" => DATA <= x"7000";
            when "00" & x"d73" => DATA <= x"5387";
            when "00" & x"d74" => DATA <= x"51c9";
            when "00" & x"d75" => DATA <= x"fff6";
            when "00" & x"d76" => DATA <= x"9487";
            when "00" & x"d77" => DATA <= x"1dbc";
            when "00" & x"d78" => DATA <= x"0020";
            when "00" & x"d79" => DATA <= x"7000";
            when "00" & x"d7a" => DATA <= x"51cf";
            when "00" & x"d7b" => DATA <= x"fff8";
            when "00" & x"d7c" => DATA <= x"201f";
            when "00" & x"d7d" => DATA <= x"221f";
            when "00" & x"d7e" => DATA <= x"2c5f";
            when "00" & x"d7f" => DATA <= x"4e75";
            when "00" & x"d80" => DATA <= x"203c";
            when "00" & x"d81" => DATA <= x"003f";
            when "00" & x"d82" => DATA <= x"2e80";
            when "00" & x"d83" => DATA <= x"003c";
            when "00" & x"d84" => DATA <= x"0002";
            when "00" & x"d85" => DATA <= x"4e75";
            when "00" & x"d86" => DATA <= x"2f03";
            when "00" & x"d87" => DATA <= x"2f00";
            when "00" & x"d88" => DATA <= x"0280";
            when "00" & x"d89" => DATA <= x"0000";
            when "00" & x"d8a" => DATA <= x"0001";
            when "00" & x"d8b" => DATA <= x"6600";
            when "00" & x"d8c" => DATA <= x"002c";
            when "00" & x"d8d" => DATA <= x"201f";
            when "00" & x"d8e" => DATA <= x"c188";
            when "00" & x"d8f" => DATA <= x"c389";
            when "00" & x"d90" => DATA <= x"2c7c";
            when "00" & x"d91" => DATA <= x"003f";
            when "00" & x"d92" => DATA <= x"39e0";
            when "00" & x"d93" => DATA <= x"3610";
            when "00" & x"d94" => DATA <= x"c66e";
            when "00" & x"d95" => DATA <= x"0002";
            when "00" & x"d96" => DATA <= x"b656";
            when "00" & x"d97" => DATA <= x"6700";
            when "00" & x"d98" => DATA <= x"000a";
            when "00" & x"d99" => DATA <= x"ddfc";
            when "00" & x"d9a" => DATA <= x"0000";
            when "00" & x"d9b" => DATA <= x"000e";
            when "00" & x"d9c" => DATA <= x"60ec";
            when "00" & x"d9d" => DATA <= x"588e";
            when "00" & x"d9e" => DATA <= x"12de";
            when "00" & x"d9f" => DATA <= x"66fc";
            when "00" & x"da0" => DATA <= x"261f";
            when "00" & x"da1" => DATA <= x"4e75";
            when "00" & x"da2" => DATA <= x"261f";
            when "00" & x"da3" => DATA <= x"203c";
            when "00" & x"da4" => DATA <= x"003f";
            when "00" & x"da5" => DATA <= x"2f0c";
            when "00" & x"da6" => DATA <= x"003c";
            when "00" & x"da7" => DATA <= x"0002";
            when "00" & x"da8" => DATA <= x"4e75";
            when "00" & x"da9" => DATA <= x"0c16";
            when "00" & x"daa" => DATA <= x"000d";
            when "00" & x"dab" => DATA <= x"6700";
            when "00" & x"dac" => DATA <= x"004c";
            when "00" & x"dad" => DATA <= x"2f0e";
            when "00" & x"dae" => DATA <= x"7010";
            when "00" & x"daf" => DATA <= x"220e";
            when "00" & x"db0" => DATA <= x"6100";
            when "00" & x"db1" => DATA <= x"f46a";
            when "00" & x"db2" => DATA <= x"6800";
            when "00" & x"db3" => DATA <= x"0010";
            when "00" & x"db4" => DATA <= x"21fc";
            when "00" & x"db5" => DATA <= x"0000";
            when "00" & x"db6" => DATA <= x"0000";
            when "00" & x"db7" => DATA <= x"0700";
            when "00" & x"db8" => DATA <= x"2c5f";
            when "00" & x"db9" => DATA <= x"6000";
            when "00" & x"dba" => DATA <= x"000a";
            when "00" & x"dbb" => DATA <= x"2c41";
            when "00" & x"dbc" => DATA <= x"21c2";
            when "00" & x"dbd" => DATA <= x"0700";
            when "00" & x"dbe" => DATA <= x"241f";
            when "00" & x"dbf" => DATA <= x"6100";
            when "00" & x"dc0" => DATA <= x"0ba0";
            when "00" & x"dc1" => DATA <= x"6500";
            when "00" & x"dc2" => DATA <= x"0020";
            when "00" & x"dc3" => DATA <= x"2a7c";
            when "00" & x"dc4" => DATA <= x"0000";
            when "00" & x"dc5" => DATA <= x"0704";
            when "00" & x"dc6" => DATA <= x"1a9e";
            when "00" & x"dc7" => DATA <= x"0c1d";
            when "00" & x"dc8" => DATA <= x"000d";
            when "00" & x"dc9" => DATA <= x"66f8";
            when "00" & x"dca" => DATA <= x"1b3c";
            when "00" & x"dcb" => DATA <= x"0000";
            when "00" & x"dcc" => DATA <= x"203c";
            when "00" & x"dcd" => DATA <= x"0000";
            when "00" & x"dce" => DATA <= x"0700";
            when "00" & x"dcf" => DATA <= x"6100";
            when "00" & x"dd0" => DATA <= x"f580";
            when "00" & x"dd1" => DATA <= x"4e75";
            when "00" & x"dd2" => DATA <= x"203c";
            when "00" & x"dd3" => DATA <= x"003f";
            when "00" & x"dd4" => DATA <= x"28f8";
            when "00" & x"dd5" => DATA <= x"6100";
            when "00" & x"dd6" => DATA <= x"ee52";
            when "00" & x"dd7" => DATA <= x"4e75";
            when "00" & x"dd8" => DATA <= x"2f0e";
            when "00" & x"dd9" => DATA <= x"6100";
            when "00" & x"dda" => DATA <= x"0b6c";
            when "00" & x"ddb" => DATA <= x"0c16";
            when "00" & x"ddc" => DATA <= x"000d";
            when "00" & x"ddd" => DATA <= x"6700";
            when "00" & x"dde" => DATA <= x"0010";
            when "00" & x"ddf" => DATA <= x"0c16";
            when "00" & x"de0" => DATA <= x"000d";
            when "00" & x"de1" => DATA <= x"6700";
            when "00" & x"de2" => DATA <= x"0016";
            when "00" & x"de3" => DATA <= x"0c1e";
            when "00" & x"de4" => DATA <= x"0020";
            when "00" & x"de5" => DATA <= x"66f2";
            when "00" & x"de6" => DATA <= x"203c";
            when "00" & x"de7" => DATA <= x"003f";
            when "00" & x"de8" => DATA <= x"2bfe";
            when "00" & x"de9" => DATA <= x"6100";
            when "00" & x"dea" => DATA <= x"ee2a";
            when "00" & x"deb" => DATA <= x"2c5f";
            when "00" & x"dec" => DATA <= x"4e75";
            when "00" & x"ded" => DATA <= x"2c5f";
            when "00" & x"dee" => DATA <= x"220e";
            when "00" & x"def" => DATA <= x"7005";
            when "00" & x"df0" => DATA <= x"6100";
            when "00" & x"df1" => DATA <= x"f0e8";
            when "00" & x"df2" => DATA <= x"b8bc";
            when "00" & x"df3" => DATA <= x"0000";
            when "00" & x"df4" => DATA <= x"8000";
            when "00" & x"df5" => DATA <= x"6600";
            when "00" & x"df6" => DATA <= x"0078";
            when "00" & x"df7" => DATA <= x"2a78";
            when "00" & x"df8" => DATA <= x"0504";
            when "00" & x"df9" => DATA <= x"dbfc";
            when "00" & x"dfa" => DATA <= x"0000";
            when "00" & x"dfb" => DATA <= x"8000";
            when "00" & x"dfc" => DATA <= x"dbfc";
            when "00" & x"dfd" => DATA <= x"0000";
            when "00" & x"dfe" => DATA <= x"0100";
            when "00" & x"dff" => DATA <= x"bbf8";
            when "00" & x"e00" => DATA <= x"0508";
            when "00" & x"e01" => DATA <= x"6300";
            when "00" & x"e02" => DATA <= x"006c";
            when "00" & x"e03" => DATA <= x"220e";
            when "00" & x"e04" => DATA <= x"243c";
            when "00" & x"e05" => DATA <= x"0000";
            when "00" & x"e06" => DATA <= x"0400";
            when "00" & x"e07" => DATA <= x"7600";
            when "00" & x"e08" => DATA <= x"203c";
            when "00" & x"e09" => DATA <= x"0000";
            when "00" & x"e0a" => DATA <= x"00ff";
            when "00" & x"e0b" => DATA <= x"6100";
            when "00" & x"e0c" => DATA <= x"f0b2";
            when "00" & x"e0d" => DATA <= x"203c";
            when "00" & x"e0e" => DATA <= x"003f";
            when "00" & x"e0f" => DATA <= x"2b5d";
            when "00" & x"e10" => DATA <= x"6100";
            when "00" & x"e11" => DATA <= x"eddc";
            when "00" & x"e12" => DATA <= x"7015";
            when "00" & x"e13" => DATA <= x"7200";
            when "00" & x"e14" => DATA <= x"6100";
            when "00" & x"e15" => DATA <= x"eea8";
            when "00" & x"e16" => DATA <= x"6100";
            when "00" & x"e17" => DATA <= x"f86c";
            when "00" & x"e18" => DATA <= x"6100";
            when "00" & x"e19" => DATA <= x"edb4";
            when "00" & x"e1a" => DATA <= x"66a0";
            when "00" & x"e1b" => DATA <= x"223c";
            when "00" & x"e1c" => DATA <= x"0000";
            when "00" & x"e1d" => DATA <= x"0600";
            when "00" & x"e1e" => DATA <= x"74ff";
            when "00" & x"e1f" => DATA <= x"203c";
            when "00" & x"e20" => DATA <= x"003f";
            when "00" & x"e21" => DATA <= x"2bca";
            when "00" & x"e22" => DATA <= x"6100";
            when "00" & x"e23" => DATA <= x"edb8";
            when "00" & x"e24" => DATA <= x"1007";
            when "00" & x"e25" => DATA <= x"0600";
            when "00" & x"e26" => DATA <= x"0030";
            when "00" & x"e27" => DATA <= x"6100";
            when "00" & x"e28" => DATA <= x"ed96";
            when "00" & x"e29" => DATA <= x"6100";
            when "00" & x"e2a" => DATA <= x"edbe";
            when "00" & x"e2b" => DATA <= x"203c";
            when "00" & x"e2c" => DATA <= x"003f";
            when "00" & x"e2d" => DATA <= x"2bdf";
            when "00" & x"e2e" => DATA <= x"6100";
            when "00" & x"e2f" => DATA <= x"eda0";
            when "00" & x"e30" => DATA <= x"6000";
            when "00" & x"e31" => DATA <= x"ff74";
            when "00" & x"e32" => DATA <= x"203c";
            when "00" & x"e33" => DATA <= x"003f";
            when "00" & x"e34" => DATA <= x"2b37";
            when "00" & x"e35" => DATA <= x"6100";
            when "00" & x"e36" => DATA <= x"ed92";
            when "00" & x"e37" => DATA <= x"4e75";
            when "00" & x"e38" => DATA <= x"203c";
            when "00" & x"e39" => DATA <= x"003f";
            when "00" & x"e3a" => DATA <= x"2b53";
            when "00" & x"e3b" => DATA <= x"6100";
            when "00" & x"e3c" => DATA <= x"ed86";
            when "00" & x"e3d" => DATA <= x"4e75";
            when "00" & x"e3e" => DATA <= x"203c";
            when "00" & x"e3f" => DATA <= x"003f";
            when "00" & x"e40" => DATA <= x"291b";
            when "00" & x"e41" => DATA <= x"6100";
            when "00" & x"e42" => DATA <= x"ed7a";
            when "00" & x"e43" => DATA <= x"4e75";
            when "00" & x"e44" => DATA <= x"7010";
            when "00" & x"e45" => DATA <= x"220e";
            when "00" & x"e46" => DATA <= x"6100";
            when "00" & x"e47" => DATA <= x"f33e";
            when "00" & x"e48" => DATA <= x"6900";
            when "00" & x"e49" => DATA <= x"0018";
            when "00" & x"e4a" => DATA <= x"6100";
            when "00" & x"e4b" => DATA <= x"0a98";
            when "00" & x"e4c" => DATA <= x"6600";
            when "00" & x"e4d" => DATA <= x"0010";
            when "00" & x"e4e" => DATA <= x"21c2";
            when "00" & x"e4f" => DATA <= x"0520";
            when "00" & x"e50" => DATA <= x"6100";
            when "00" & x"e51" => DATA <= x"eee2";
            when "00" & x"e52" => DATA <= x"023c";
            when "00" & x"e53" => DATA <= x"00fe";
            when "00" & x"e54" => DATA <= x"4e75";
            when "00" & x"e55" => DATA <= x"203c";
            when "00" & x"e56" => DATA <= x"003f";
            when "00" & x"e57" => DATA <= x"2931";
            when "00" & x"e58" => DATA <= x"6100";
            when "00" & x"e59" => DATA <= x"ed4c";
            when "00" & x"e5a" => DATA <= x"4e75";
            when "00" & x"e5b" => DATA <= x"2f0e";
            when "00" & x"e5c" => DATA <= x"0c16";
            when "00" & x"e5d" => DATA <= x"000d";
            when "00" & x"e5e" => DATA <= x"6600";
            when "00" & x"e5f" => DATA <= x"001a";
            when "00" & x"e60" => DATA <= x"203c";
            when "00" & x"e61" => DATA <= x"003f";
            when "00" & x"e62" => DATA <= x"2838";
            when "00" & x"e63" => DATA <= x"6100";
            when "00" & x"e64" => DATA <= x"ed36";
            when "00" & x"e65" => DATA <= x"203c";
            when "00" & x"e66" => DATA <= x"003f";
            when "00" & x"e67" => DATA <= x"2859";
            when "00" & x"e68" => DATA <= x"6100";
            when "00" & x"e69" => DATA <= x"ed2c";
            when "00" & x"e6a" => DATA <= x"6000";
            when "00" & x"e6b" => DATA <= x"00ca";
            when "00" & x"e6c" => DATA <= x"0216";
            when "00" & x"e6d" => DATA <= x"00df";
            when "00" & x"e6e" => DATA <= x"0c1e";
            when "00" & x"e6f" => DATA <= x"0054";
            when "00" & x"e70" => DATA <= x"6600";
            when "00" & x"e71" => DATA <= x"0042";
            when "00" & x"e72" => DATA <= x"0216";
            when "00" & x"e73" => DATA <= x"00df";
            when "00" & x"e74" => DATA <= x"0c1e";
            when "00" & x"e75" => DATA <= x"0055";
            when "00" & x"e76" => DATA <= x"6600";
            when "00" & x"e77" => DATA <= x"00b2";
            when "00" & x"e78" => DATA <= x"0216";
            when "00" & x"e79" => DATA <= x"00df";
            when "00" & x"e7a" => DATA <= x"0c1e";
            when "00" & x"e7b" => DATA <= x"0042";
            when "00" & x"e7c" => DATA <= x"6600";
            when "00" & x"e7d" => DATA <= x"00a6";
            when "00" & x"e7e" => DATA <= x"0216";
            when "00" & x"e7f" => DATA <= x"00df";
            when "00" & x"e80" => DATA <= x"0c1e";
            when "00" & x"e81" => DATA <= x"0045";
            when "00" & x"e82" => DATA <= x"6600";
            when "00" & x"e83" => DATA <= x"009a";
            when "00" & x"e84" => DATA <= x"0c16";
            when "00" & x"e85" => DATA <= x"000d";
            when "00" & x"e86" => DATA <= x"6600";
            when "00" & x"e87" => DATA <= x"0092";
            when "00" & x"e88" => DATA <= x"203c";
            when "00" & x"e89" => DATA <= x"003f";
            when "00" & x"e8a" => DATA <= x"2838";
            when "00" & x"e8b" => DATA <= x"6100";
            when "00" & x"e8c" => DATA <= x"ece6";
            when "00" & x"e8d" => DATA <= x"203c";
            when "00" & x"e8e" => DATA <= x"003f";
            when "00" & x"e8f" => DATA <= x"286b";
            when "00" & x"e90" => DATA <= x"6100";
            when "00" & x"e91" => DATA <= x"ecdc";
            when "00" & x"e92" => DATA <= x"0226";
            when "00" & x"e93" => DATA <= x"00df";
            when "00" & x"e94" => DATA <= x"0c1e";
            when "00" & x"e95" => DATA <= x"0053";
            when "00" & x"e96" => DATA <= x"6600";
            when "00" & x"e97" => DATA <= x"0072";
            when "00" & x"e98" => DATA <= x"0216";
            when "00" & x"e99" => DATA <= x"00df";
            when "00" & x"e9a" => DATA <= x"0c1e";
            when "00" & x"e9b" => DATA <= x"0057";
            when "00" & x"e9c" => DATA <= x"6600";
            when "00" & x"e9d" => DATA <= x"0066";
            when "00" & x"e9e" => DATA <= x"0216";
            when "00" & x"e9f" => DATA <= x"00df";
            when "00" & x"ea0" => DATA <= x"0c1e";
            when "00" & x"ea1" => DATA <= x"0049";
            when "00" & x"ea2" => DATA <= x"6600";
            when "00" & x"ea3" => DATA <= x"005a";
            when "00" & x"ea4" => DATA <= x"0c16";
            when "00" & x"ea5" => DATA <= x"000d";
            when "00" & x"ea6" => DATA <= x"6600";
            when "00" & x"ea7" => DATA <= x"0052";
            when "00" & x"ea8" => DATA <= x"203c";
            when "00" & x"ea9" => DATA <= x"003f";
            when "00" & x"eaa" => DATA <= x"2838";
            when "00" & x"eab" => DATA <= x"6100";
            when "00" & x"eac" => DATA <= x"eca6";
            when "00" & x"ead" => DATA <= x"4df9";
            when "00" & x"eae" => DATA <= x"003f";
            when "00" & x"eaf" => DATA <= x"2f50";
            when "00" & x"eb0" => DATA <= x"103c";
            when "00" & x"eb1" => DATA <= x"0020";
            when "00" & x"eb2" => DATA <= x"6100";
            when "00" & x"eb3" => DATA <= x"ec80";
            when "00" & x"eb4" => DATA <= x"6100";
            when "00" & x"eb5" => DATA <= x"ec7c";
            when "00" & x"eb6" => DATA <= x"6100";
            when "00" & x"eb7" => DATA <= x"ec78";
            when "00" & x"eb8" => DATA <= x"201e";
            when "00" & x"eb9" => DATA <= x"201e";
            when "00" & x"eba" => DATA <= x"0c80";
            when "00" & x"ebb" => DATA <= x"ffff";
            when "00" & x"ebc" => DATA <= x"ffff";
            when "00" & x"ebd" => DATA <= x"6700";
            when "00" & x"ebe" => DATA <= x"0024";
            when "00" & x"ebf" => DATA <= x"200e";
            when "00" & x"ec0" => DATA <= x"6100";
            when "00" & x"ec1" => DATA <= x"ec7c";
            when "00" & x"ec2" => DATA <= x"2c40";
            when "00" & x"ec3" => DATA <= x"0c26";
            when "00" & x"ec4" => DATA <= x"0000";
            when "00" & x"ec5" => DATA <= x"6100";
            when "00" & x"ec6" => DATA <= x"ec86";
            when "00" & x"ec7" => DATA <= x"0c1e";
            when "00" & x"ec8" => DATA <= x"00ff";
            when "00" & x"ec9" => DATA <= x"6700";
            when "00" & x"eca" => DATA <= x"000c";
            when "00" & x"ecb" => DATA <= x"200e";
            when "00" & x"ecc" => DATA <= x"0200";
            when "00" & x"ecd" => DATA <= x"0003";
            when "00" & x"ece" => DATA <= x"66f0";
            when "00" & x"ecf" => DATA <= x"60c0";
            when "00" & x"ed0" => DATA <= x"2f01";
            when "00" & x"ed1" => DATA <= x"7209";
            when "00" & x"ed2" => DATA <= x"6100";
            when "00" & x"ed3" => DATA <= x"f3aa";
            when "00" & x"ed4" => DATA <= x"221f";
            when "00" & x"ed5" => DATA <= x"2c5f";
            when "00" & x"ed6" => DATA <= x"003c";
            when "00" & x"ed7" => DATA <= x"0001";
            when "00" & x"ed8" => DATA <= x"4e75";
            when "00" & x"ed9" => DATA <= x"0c16";
            when "00" & x"eda" => DATA <= x"000d";
            when "00" & x"edb" => DATA <= x"6600";
            when "00" & x"edc" => DATA <= x"06b8";
            when "00" & x"edd" => DATA <= x"203c";
            when "00" & x"ede" => DATA <= x"003f";
            when "00" & x"edf" => DATA <= x"299f";
            when "00" & x"ee0" => DATA <= x"6100";
            when "00" & x"ee1" => DATA <= x"ec3c";
            when "00" & x"ee2" => DATA <= x"6100";
            when "00" & x"ee3" => DATA <= x"ec4c";
            when "00" & x"ee4" => DATA <= x"103c";
            when "00" & x"ee5" => DATA <= x"003a";
            when "00" & x"ee6" => DATA <= x"6100";
            when "00" & x"ee7" => DATA <= x"ec18";
            when "00" & x"ee8" => DATA <= x"203c";
            when "00" & x"ee9" => DATA <= x"0000";
            when "00" & x"eea" => DATA <= x"0600";
            when "00" & x"eeb" => DATA <= x"123c";
            when "00" & x"eec" => DATA <= x"00ff";
            when "00" & x"eed" => DATA <= x"143c";
            when "00" & x"eee" => DATA <= x"0020";
            when "00" & x"eef" => DATA <= x"163c";
            when "00" & x"ef0" => DATA <= x"00ff";
            when "00" & x"ef1" => DATA <= x"207c";
            when "00" & x"ef2" => DATA <= x"0000";
            when "00" & x"ef3" => DATA <= x"007d";
            when "00" & x"ef4" => DATA <= x"4e4c";
            when "00" & x"ef5" => DATA <= x"6500";
            when "00" & x"ef6" => DATA <= x"00b8";
            when "00" & x"ef7" => DATA <= x"2c7c";
            when "00" & x"ef8" => DATA <= x"0000";
            when "00" & x"ef9" => DATA <= x"0600";
            when "00" & x"efa" => DATA <= x"101e";
            when "00" & x"efb" => DATA <= x"b03c";
            when "00" & x"efc" => DATA <= x"003f";
            when "00" & x"efd" => DATA <= x"6700";
            when "00" & x"efe" => DATA <= x"02c8";
            when "00" & x"eff" => DATA <= x"b03c";
            when "00" & x"f00" => DATA <= x"002a";
            when "00" & x"f01" => DATA <= x"6700";
            when "00" & x"f02" => DATA <= x"03b2";
            when "00" & x"f03" => DATA <= x"0200";
            when "00" & x"f04" => DATA <= x"00df";
            when "00" & x"f05" => DATA <= x"b03c";
            when "00" & x"f06" => DATA <= x"0042";
            when "00" & x"f07" => DATA <= x"6700";
            when "00" & x"f08" => DATA <= x"009e";
            when "00" & x"f09" => DATA <= x"b03c";
            when "00" & x"f0a" => DATA <= x"0044";
            when "00" & x"f0b" => DATA <= x"6700";
            when "00" & x"f0c" => DATA <= x"0060";
            when "00" & x"f0d" => DATA <= x"b03c";
            when "00" & x"f0e" => DATA <= x"0045";
            when "00" & x"f0f" => DATA <= x"6700";
            when "00" & x"f10" => DATA <= x"00f2";
            when "00" & x"f11" => DATA <= x"b03c";
            when "00" & x"f12" => DATA <= x"0046";
            when "00" & x"f13" => DATA <= x"6700";
            when "00" & x"f14" => DATA <= x"01a0";
            when "00" & x"f15" => DATA <= x"b03c";
            when "00" & x"f16" => DATA <= x"0047";
            when "00" & x"f17" => DATA <= x"6700";
            when "00" & x"f18" => DATA <= x"01d2";
            when "00" & x"f19" => DATA <= x"b03c";
            when "00" & x"f1a" => DATA <= x"0048";
            when "00" & x"f1b" => DATA <= x"6700";
            when "00" & x"f1c" => DATA <= x"01e6";
            when "00" & x"f1d" => DATA <= x"b03c";
            when "00" & x"f1e" => DATA <= x"004d";
            when "00" & x"f1f" => DATA <= x"6700";
            when "00" & x"f20" => DATA <= x"0292";
            when "00" & x"f21" => DATA <= x"b03c";
            when "00" & x"f22" => DATA <= x"0051";
            when "00" & x"f23" => DATA <= x"6700";
            when "00" & x"f24" => DATA <= x"02c0";
            when "00" & x"f25" => DATA <= x"b03c";
            when "00" & x"f26" => DATA <= x"0052";
            when "00" & x"f27" => DATA <= x"6700";
            when "00" & x"f28" => DATA <= x"02be";
            when "00" & x"f29" => DATA <= x"b03c";
            when "00" & x"f2a" => DATA <= x"0053";
            when "00" & x"f2b" => DATA <= x"6700";
            when "00" & x"f2c" => DATA <= x"0012";
            when "00" & x"f2d" => DATA <= x"b03c";
            when "00" & x"f2e" => DATA <= x"0054";
            when "00" & x"f2f" => DATA <= x"6700";
            when "00" & x"f30" => DATA <= x"000a";
            when "00" & x"f31" => DATA <= x"b03c";
            when "00" & x"f32" => DATA <= x"0056";
            when "00" & x"f33" => DATA <= x"6700";
            when "00" & x"f34" => DATA <= x"0358";
            when "00" & x"f35" => DATA <= x"203c";
            when "00" & x"f36" => DATA <= x"003f";
            when "00" & x"f37" => DATA <= x"2b03";
            when "00" & x"f38" => DATA <= x"6100";
            when "00" & x"f39" => DATA <= x"eb8c";
            when "00" & x"f3a" => DATA <= x"6000";
            when "00" & x"f3b" => DATA <= x"ff4e";
            when "00" & x"f3c" => DATA <= x"6100";
            when "00" & x"f3d" => DATA <= x"08a6";
            when "00" & x"f3e" => DATA <= x"7010";
            when "00" & x"f3f" => DATA <= x"220e";
            when "00" & x"f40" => DATA <= x"6100";
            when "00" & x"f41" => DATA <= x"f14a";
            when "00" & x"f42" => DATA <= x"6900";
            when "00" & x"f43" => DATA <= x"023e";
            when "00" & x"f44" => DATA <= x"2c41";
            when "00" & x"f45" => DATA <= x"2002";
            when "00" & x"f46" => DATA <= x"223c";
            when "00" & x"f47" => DATA <= x"0000";
            when "00" & x"f48" => DATA <= x"0600";
            when "00" & x"f49" => DATA <= x"6100";
            when "00" & x"f4a" => DATA <= x"fc78";
            when "00" & x"f4b" => DATA <= x"2001";
            when "00" & x"f4c" => DATA <= x"6100";
            when "00" & x"f4d" => DATA <= x"eb64";
            when "00" & x"f4e" => DATA <= x"6100";
            when "00" & x"f4f" => DATA <= x"eb74";
            when "00" & x"f50" => DATA <= x"6000";
            when "00" & x"f51" => DATA <= x"ff22";
            when "00" & x"f52" => DATA <= x"707e";
            when "00" & x"f53" => DATA <= x"6100";
            when "00" & x"f54" => DATA <= x"ec2a";
            when "00" & x"f55" => DATA <= x"6000";
            when "00" & x"f56" => DATA <= x"ff18";
            when "00" & x"f57" => DATA <= x"6100";
            when "00" & x"f58" => DATA <= x"0870";
            when "00" & x"f59" => DATA <= x"7010";
            when "00" & x"f5a" => DATA <= x"220e";
            when "00" & x"f5b" => DATA <= x"6100";
            when "00" & x"f5c" => DATA <= x"f114";
            when "00" & x"f5d" => DATA <= x"6900";
            when "00" & x"f5e" => DATA <= x"0208";
            when "00" & x"f5f" => DATA <= x"2842";
            when "00" & x"f60" => DATA <= x"6100";
            when "00" & x"f61" => DATA <= x"086c";
            when "00" & x"f62" => DATA <= x"7010";
            when "00" & x"f63" => DATA <= x"6100";
            when "00" & x"f64" => DATA <= x"f104";
            when "00" & x"f65" => DATA <= x"6900";
            when "00" & x"f66" => DATA <= x"01f8";
            when "00" & x"f67" => DATA <= x"2a42";
            when "00" & x"f68" => DATA <= x"6100";
            when "00" & x"f69" => DATA <= x"085c";
            when "00" & x"f6a" => DATA <= x"7010";
            when "00" & x"f6b" => DATA <= x"6100";
            when "00" & x"f6c" => DATA <= x"f0f4";
            when "00" & x"f6d" => DATA <= x"6900";
            when "00" & x"f6e" => DATA <= x"01e8";
            when "00" & x"f6f" => DATA <= x"2c41";
            when "00" & x"f70" => DATA <= x"1e02";
            when "00" & x"f71" => DATA <= x"be1c";
            when "00" & x"f72" => DATA <= x"6600";
            when "00" & x"f73" => DATA <= x"0024";
            when "00" & x"f74" => DATA <= x"200c";
            when "00" & x"f75" => DATA <= x"223c";
            when "00" & x"f76" => DATA <= x"0000";
            when "00" & x"f77" => DATA <= x"0600";
            when "00" & x"f78" => DATA <= x"243c";
            when "00" & x"f79" => DATA <= x"0000";
            when "00" & x"f7a" => DATA <= x"00ff";
            when "00" & x"f7b" => DATA <= x"6100";
            when "00" & x"f7c" => DATA <= x"f7ee";
            when "00" & x"f7d" => DATA <= x"21fc";
            when "00" & x"f7e" => DATA <= x"2020";
            when "00" & x"f7f" => DATA <= x"0000";
            when "00" & x"f80" => DATA <= x"0608";
            when "00" & x"f81" => DATA <= x"303c";
            when "00" & x"f82" => DATA <= x"0600";
            when "00" & x"f83" => DATA <= x"6100";
            when "00" & x"f84" => DATA <= x"eaf6";
            when "00" & x"f85" => DATA <= x"bbcc";
            when "00" & x"f86" => DATA <= x"64d4";
            when "00" & x"f87" => DATA <= x"6000";
            when "00" & x"f88" => DATA <= x"feb4";
            when "00" & x"f89" => DATA <= x"6100";
            when "00" & x"f8a" => DATA <= x"080c";
            when "00" & x"f8b" => DATA <= x"7010";
            when "00" & x"f8c" => DATA <= x"220e";
            when "00" & x"f8d" => DATA <= x"6100";
            when "00" & x"f8e" => DATA <= x"f0b0";
            when "00" & x"f8f" => DATA <= x"6900";
            when "00" & x"f90" => DATA <= x"01a4";
            when "00" & x"f91" => DATA <= x"2842";
            when "00" & x"f92" => DATA <= x"11fc";
            when "00" & x"f93" => DATA <= x"0020";
            when "00" & x"f94" => DATA <= x"0609";
            when "00" & x"f95" => DATA <= x"11fc";
            when "00" & x"f96" => DATA <= x"0020";
            when "00" & x"f97" => DATA <= x"060d";
            when "00" & x"f98" => DATA <= x"11fc";
            when "00" & x"f99" => DATA <= x"0028";
            when "00" & x"f9a" => DATA <= x"060e";
            when "00" & x"f9b" => DATA <= x"21fc";
            when "00" & x"f9c" => DATA <= x"2920";
            when "00" & x"f9d" => DATA <= x"2000";
            when "00" & x"f9e" => DATA <= x"0610";
            when "00" & x"f9f" => DATA <= x"200c";
            when "00" & x"fa0" => DATA <= x"223c";
            when "00" & x"fa1" => DATA <= x"0000";
            when "00" & x"fa2" => DATA <= x"0600";
            when "00" & x"fa3" => DATA <= x"243c";
            when "00" & x"fa4" => DATA <= x"0000";
            when "00" & x"fa5" => DATA <= x"00ff";
            when "00" & x"fa6" => DATA <= x"6100";
            when "00" & x"fa7" => DATA <= x"f798";
            when "00" & x"fa8" => DATA <= x"11fc";
            when "00" & x"fa9" => DATA <= x"0020";
            when "00" & x"faa" => DATA <= x"0608";
            when "00" & x"fab" => DATA <= x"5441";
            when "00" & x"fac" => DATA <= x"1014";
            when "00" & x"fad" => DATA <= x"243c";
            when "00" & x"fae" => DATA <= x"0000";
            when "00" & x"faf" => DATA <= x"00ff";
            when "00" & x"fb0" => DATA <= x"6100";
            when "00" & x"fb1" => DATA <= x"f72e";
            when "00" & x"fb2" => DATA <= x"2a41";
            when "00" & x"fb3" => DATA <= x"1afc";
            when "00" & x"fb4" => DATA <= x"0020";
            when "00" & x"fb5" => DATA <= x"2c4c";
            when "00" & x"fb6" => DATA <= x"6100";
            when "00" & x"fb7" => DATA <= x"084c";
            when "00" & x"fb8" => DATA <= x"11c0";
            when "00" & x"fb9" => DATA <= x"060f";
            when "00" & x"fba" => DATA <= x"203c";
            when "00" & x"fbb" => DATA <= x"0000";
            when "00" & x"fbc" => DATA <= x"0600";
            when "00" & x"fbd" => DATA <= x"6100";
            when "00" & x"fbe" => DATA <= x"ea82";
            when "00" & x"fbf" => DATA <= x"203c";
            when "00" & x"fc0" => DATA <= x"0000";
            when "00" & x"fc1" => DATA <= x"0680";
            when "00" & x"fc2" => DATA <= x"123c";
            when "00" & x"fc3" => DATA <= x"0002";
            when "00" & x"fc4" => DATA <= x"143c";
            when "00" & x"fc5" => DATA <= x"0020";
            when "00" & x"fc6" => DATA <= x"163c";
            when "00" & x"fc7" => DATA <= x"0046";
            when "00" & x"fc8" => DATA <= x"207c";
            when "00" & x"fc9" => DATA <= x"0000";
            when "00" & x"fca" => DATA <= x"007d";
            when "00" & x"fcb" => DATA <= x"4e4c";
            when "00" & x"fcc" => DATA <= x"6500";
            when "00" & x"fcd" => DATA <= x"0024";
            when "00" & x"fce" => DATA <= x"0c38";
            when "00" & x"fcf" => DATA <= x"000d";
            when "00" & x"fd0" => DATA <= x"0680";
            when "00" & x"fd1" => DATA <= x"6600";
            when "00" & x"fd2" => DATA <= x"0006";
            when "00" & x"fd3" => DATA <= x"524c";
            when "00" & x"fd4" => DATA <= x"6094";
            when "00" & x"fd5" => DATA <= x"2c7c";
            when "00" & x"fd6" => DATA <= x"0000";
            when "00" & x"fd7" => DATA <= x"0680";
            when "00" & x"fd8" => DATA <= x"7010";
            when "00" & x"fd9" => DATA <= x"220e";
            when "00" & x"fda" => DATA <= x"6100";
            when "00" & x"fdb" => DATA <= x"f016";
            when "00" & x"fdc" => DATA <= x"6984";
            when "00" & x"fdd" => DATA <= x"18c2";
            when "00" & x"fde" => DATA <= x"6080";
            when "00" & x"fdf" => DATA <= x"707e";
            when "00" & x"fe0" => DATA <= x"6100";
            when "00" & x"fe1" => DATA <= x"eb10";
            when "00" & x"fe2" => DATA <= x"6000";
            when "00" & x"fe3" => DATA <= x"fdfe";
            when "00" & x"fe4" => DATA <= x"220e";
            when "00" & x"fe5" => DATA <= x"6100";
            when "00" & x"fe6" => DATA <= x"0762";
            when "00" & x"fe7" => DATA <= x"7010";
            when "00" & x"fe8" => DATA <= x"6100";
            when "00" & x"fe9" => DATA <= x"effa";
            when "00" & x"fea" => DATA <= x"6900";
            when "00" & x"feb" => DATA <= x"00ee";
            when "00" & x"fec" => DATA <= x"2842";
            when "00" & x"fed" => DATA <= x"6100";
            when "00" & x"fee" => DATA <= x"0752";
            when "00" & x"fef" => DATA <= x"7010";
            when "00" & x"ff0" => DATA <= x"6100";
            when "00" & x"ff1" => DATA <= x"efea";
            when "00" & x"ff2" => DATA <= x"6900";
            when "00" & x"ff3" => DATA <= x"00de";
            when "00" & x"ff4" => DATA <= x"2a42";
            when "00" & x"ff5" => DATA <= x"6100";
            when "00" & x"ff6" => DATA <= x"0742";
            when "00" & x"ff7" => DATA <= x"7010";
            when "00" & x"ff8" => DATA <= x"6100";
            when "00" & x"ff9" => DATA <= x"efda";
            when "00" & x"ffa" => DATA <= x"6900";
            when "00" & x"ffb" => DATA <= x"00ce";
            when "00" & x"ffc" => DATA <= x"18c2";
            when "00" & x"ffd" => DATA <= x"bbcc";
            when "00" & x"ffe" => DATA <= x"64fa";
            when "00" & x"fff" => DATA <= x"6000";
            when "01" & x"000" => DATA <= x"fdc4";
            when "01" & x"001" => DATA <= x"6100";
            when "01" & x"002" => DATA <= x"071c";
            when "01" & x"003" => DATA <= x"6700";
            when "01" & x"004" => DATA <= x"00bc";
            when "01" & x"005" => DATA <= x"7010";
            when "01" & x"006" => DATA <= x"220e";
            when "01" & x"007" => DATA <= x"6100";
            when "01" & x"008" => DATA <= x"efbc";
            when "01" & x"009" => DATA <= x"6900";
            when "01" & x"00a" => DATA <= x"00b0";
            when "01" & x"00b" => DATA <= x"2c42";
            when "01" & x"00c" => DATA <= x"4e96";
            when "01" & x"00d" => DATA <= x"6000";
            when "01" & x"00e" => DATA <= x"fda8";
            when "01" & x"00f" => DATA <= x"6100";
            when "01" & x"010" => DATA <= x"0700";
            when "01" & x"011" => DATA <= x"0c16";
            when "01" & x"012" => DATA <= x"000d";
            when "01" & x"013" => DATA <= x"6600";
            when "01" & x"014" => DATA <= x"0008";
            when "01" & x"015" => DATA <= x"4282";
            when "01" & x"016" => DATA <= x"6000";
            when "01" & x"017" => DATA <= x"0016";
            when "01" & x"018" => DATA <= x"7010";
            when "01" & x"019" => DATA <= x"220e";
            when "01" & x"01a" => DATA <= x"6100";
            when "01" & x"01b" => DATA <= x"ef96";
            when "01" & x"01c" => DATA <= x"6900";
            when "01" & x"01d" => DATA <= x"008a";
            when "01" & x"01e" => DATA <= x"6100";
            when "01" & x"01f" => DATA <= x"06f0";
            when "01" & x"020" => DATA <= x"6600";
            when "01" & x"021" => DATA <= x"0082";
            when "01" & x"022" => DATA <= x"0282";
            when "01" & x"023" => DATA <= x"ffff";
            when "01" & x"024" => DATA <= x"fffc";
            when "01" & x"025" => DATA <= x"2c42";
            when "01" & x"026" => DATA <= x"103c";
            when "01" & x"027" => DATA <= x"000e";
            when "01" & x"028" => DATA <= x"6100";
            when "01" & x"029" => DATA <= x"e994";
            when "01" & x"02a" => DATA <= x"200e";
            when "01" & x"02b" => DATA <= x"223c";
            when "01" & x"02c" => DATA <= x"0000";
            when "01" & x"02d" => DATA <= x"0600";
            when "01" & x"02e" => DATA <= x"243c";
            when "01" & x"02f" => DATA <= x"0000";
            when "01" & x"030" => DATA <= x"00ff";
            when "01" & x"031" => DATA <= x"6100";
            when "01" & x"032" => DATA <= x"f682";
            when "01" & x"033" => DATA <= x"31fc";
            when "01" & x"034" => DATA <= x"2020";
            when "01" & x"035" => DATA <= x"0608";
            when "01" & x"036" => DATA <= x"5441";
            when "01" & x"037" => DATA <= x"760f";
            when "01" & x"038" => DATA <= x"287c";
            when "01" & x"039" => DATA <= x"0000";
            when "01" & x"03a" => DATA <= x"063b";
            when "01" & x"03b" => DATA <= x"11fc";
            when "01" & x"03c" => DATA <= x"0020";
            when "01" & x"03d" => DATA <= x"063a";
            when "01" & x"03e" => DATA <= x"11fc";
            when "01" & x"03f" => DATA <= x"0000";
            when "01" & x"040" => DATA <= x"064b";
            when "01" & x"041" => DATA <= x"1016";
            when "01" & x"042" => DATA <= x"243c";
            when "01" & x"043" => DATA <= x"0000";
            when "01" & x"044" => DATA <= x"00ff";
            when "01" & x"045" => DATA <= x"6100";
            when "01" & x"046" => DATA <= x"f604";
            when "01" & x"047" => DATA <= x"2a41";
            when "01" & x"048" => DATA <= x"1abc";
            when "01" & x"049" => DATA <= x"0020";
            when "01" & x"04a" => DATA <= x"5241";
            when "01" & x"04b" => DATA <= x"6100";
            when "01" & x"04c" => DATA <= x"0722";
            when "01" & x"04d" => DATA <= x"18c0";
            when "01" & x"04e" => DATA <= x"51cb";
            when "01" & x"04f" => DATA <= x"ffe4";
            when "01" & x"050" => DATA <= x"303c";
            when "01" & x"051" => DATA <= x"0600";
            when "01" & x"052" => DATA <= x"6100";
            when "01" & x"053" => DATA <= x"e958";
            when "01" & x"054" => DATA <= x"6100";
            when "01" & x"055" => DATA <= x"e968";
            when "01" & x"056" => DATA <= x"6100";
            when "01" & x"057" => DATA <= x"f078";
            when "01" & x"058" => DATA <= x"64a2";
            when "01" & x"059" => DATA <= x"707e";
            when "01" & x"05a" => DATA <= x"6100";
            when "01" & x"05b" => DATA <= x"ea1c";
            when "01" & x"05c" => DATA <= x"103c";
            when "01" & x"05d" => DATA <= x"000f";
            when "01" & x"05e" => DATA <= x"6100";
            when "01" & x"05f" => DATA <= x"e928";
            when "01" & x"060" => DATA <= x"6000";
            when "01" & x"061" => DATA <= x"fd02";
            when "01" & x"062" => DATA <= x"203c";
            when "01" & x"063" => DATA <= x"003f";
            when "01" & x"064" => DATA <= x"29ae";
            when "01" & x"065" => DATA <= x"6100";
            when "01" & x"066" => DATA <= x"e932";
            when "01" & x"067" => DATA <= x"6000";
            when "01" & x"068" => DATA <= x"fcf4";
            when "01" & x"069" => DATA <= x"6100";
            when "01" & x"06a" => DATA <= x"064c";
            when "01" & x"06b" => DATA <= x"7010";
            when "01" & x"06c" => DATA <= x"220e";
            when "01" & x"06d" => DATA <= x"6100";
            when "01" & x"06e" => DATA <= x"eef0";
            when "01" & x"06f" => DATA <= x"69e4";
            when "01" & x"070" => DATA <= x"2842";
            when "01" & x"071" => DATA <= x"6100";
            when "01" & x"072" => DATA <= x"064a";
            when "01" & x"073" => DATA <= x"7010";
            when "01" & x"074" => DATA <= x"6100";
            when "01" & x"075" => DATA <= x"eee2";
            when "01" & x"076" => DATA <= x"69d6";
            when "01" & x"077" => DATA <= x"2a42";
            when "01" & x"078" => DATA <= x"6100";
            when "01" & x"079" => DATA <= x"063c";
            when "01" & x"07a" => DATA <= x"7010";
            when "01" & x"07b" => DATA <= x"6100";
            when "01" & x"07c" => DATA <= x"eed4";
            when "01" & x"07d" => DATA <= x"69c8";
            when "01" & x"07e" => DATA <= x"5382";
            when "01" & x"07f" => DATA <= x"1adc";
            when "01" & x"080" => DATA <= x"51ca";
            when "01" & x"081" => DATA <= x"fffc";
            when "01" & x"082" => DATA <= x"6000";
            when "01" & x"083" => DATA <= x"fcbe";
            when "01" & x"084" => DATA <= x"6100";
            when "01" & x"085" => DATA <= x"e908";
            when "01" & x"086" => DATA <= x"4e75";
            when "01" & x"087" => DATA <= x"6100";
            when "01" & x"088" => DATA <= x"0610";
            when "01" & x"089" => DATA <= x"2f0d";
            when "01" & x"08a" => DATA <= x"2f02";
            when "01" & x"08b" => DATA <= x"2f01";
            when "01" & x"08c" => DATA <= x"2f00";
            when "01" & x"08d" => DATA <= x"4280";
            when "01" & x"08e" => DATA <= x"101e";
            when "01" & x"08f" => DATA <= x"0200";
            when "01" & x"090" => DATA <= x"00df";
            when "01" & x"091" => DATA <= x"0c00";
            when "01" & x"092" => DATA <= x"0041";
            when "01" & x"093" => DATA <= x"6700";
            when "01" & x"094" => DATA <= x"0008";
            when "01" & x"095" => DATA <= x"0c00";
            when "01" & x"096" => DATA <= x"0044";
            when "01" & x"097" => DATA <= x"6694";
            when "01" & x"098" => DATA <= x"0200";
            when "01" & x"099" => DATA <= x"00be";
            when "01" & x"09a" => DATA <= x"e380";
            when "01" & x"09b" => DATA <= x"1400";
            when "01" & x"09c" => DATA <= x"101e";
            when "01" & x"09d" => DATA <= x"0c00";
            when "01" & x"09e" => DATA <= x"0030";
            when "01" & x"09f" => DATA <= x"6584";
            when "01" & x"0a0" => DATA <= x"0c00";
            when "01" & x"0a1" => DATA <= x"0037";
            when "01" & x"0a2" => DATA <= x"6200";
            when "01" & x"0a3" => DATA <= x"ff7e";
            when "01" & x"0a4" => DATA <= x"0400";
            when "01" & x"0a5" => DATA <= x"0030";
            when "01" & x"0a6" => DATA <= x"d002";
            when "01" & x"0a7" => DATA <= x"e580";
            when "01" & x"0a8" => DATA <= x"2a7c";
            when "01" & x"0a9" => DATA <= x"003f";
            when "01" & x"0aa" => DATA <= x"2176";
            when "01" & x"0ab" => DATA <= x"dbc0";
            when "01" & x"0ac" => DATA <= x"6100";
            when "01" & x"0ad" => DATA <= x"05c6";
            when "01" & x"0ae" => DATA <= x"7010";
            when "01" & x"0af" => DATA <= x"220e";
            when "01" & x"0b0" => DATA <= x"6100";
            when "01" & x"0b1" => DATA <= x"ee6a";
            when "01" & x"0b2" => DATA <= x"6900";
            when "01" & x"0b3" => DATA <= x"ff5e";
            when "01" & x"0b4" => DATA <= x"4ed5";
            when "01" & x"0b5" => DATA <= x"201f";
            when "01" & x"0b6" => DATA <= x"221f";
            when "01" & x"0b7" => DATA <= x"241f";
            when "01" & x"0b8" => DATA <= x"2a5f";
            when "01" & x"0b9" => DATA <= x"6000";
            when "01" & x"0ba" => DATA <= x"fc50";
            when "01" & x"0bb" => DATA <= x"2042";
            when "01" & x"0bc" => DATA <= x"60f0";
            when "01" & x"0bd" => DATA <= x"2242";
            when "01" & x"0be" => DATA <= x"60ec";
            when "01" & x"0bf" => DATA <= x"2442";
            when "01" & x"0c0" => DATA <= x"60e8";
            when "01" & x"0c1" => DATA <= x"2642";
            when "01" & x"0c2" => DATA <= x"60e4";
            when "01" & x"0c3" => DATA <= x"2842";
            when "01" & x"0c4" => DATA <= x"60e0";
            when "01" & x"0c5" => DATA <= x"2a42";
            when "01" & x"0c6" => DATA <= x"60dc";
            when "01" & x"0c7" => DATA <= x"2c42";
            when "01" & x"0c8" => DATA <= x"60d8";
            when "01" & x"0c9" => DATA <= x"2e42";
            when "01" & x"0ca" => DATA <= x"60d4";
            when "01" & x"0cb" => DATA <= x"2002";
            when "01" & x"0cc" => DATA <= x"60d0";
            when "01" & x"0cd" => DATA <= x"2202";
            when "01" & x"0ce" => DATA <= x"60cc";
            when "01" & x"0cf" => DATA <= x"4e71";
            when "01" & x"0d0" => DATA <= x"60c8";
            when "01" & x"0d1" => DATA <= x"2602";
            when "01" & x"0d2" => DATA <= x"60c4";
            when "01" & x"0d3" => DATA <= x"2802";
            when "01" & x"0d4" => DATA <= x"60c0";
            when "01" & x"0d5" => DATA <= x"2a02";
            when "01" & x"0d6" => DATA <= x"60bc";
            when "01" & x"0d7" => DATA <= x"2c02";
            when "01" & x"0d8" => DATA <= x"60b8";
            when "01" & x"0d9" => DATA <= x"2e02";
            when "01" & x"0da" => DATA <= x"60b4";
            when "01" & x"0db" => DATA <= x"200e";
            when "01" & x"0dc" => DATA <= x"6100";
            when "01" & x"0dd" => DATA <= x"e876";
            when "01" & x"0de" => DATA <= x"6000";
            when "01" & x"0df" => DATA <= x"fc06";
            when "01" & x"0e0" => DATA <= x"103c";
            when "01" & x"0e1" => DATA <= x"0020";
            when "01" & x"0e2" => DATA <= x"323c";
            when "01" & x"0e3" => DATA <= x"0032";
            when "01" & x"0e4" => DATA <= x"6100";
            when "01" & x"0e5" => DATA <= x"e81c";
            when "01" & x"0e6" => DATA <= x"51c9";
            when "01" & x"0e7" => DATA <= x"fffa";
            when "01" & x"0e8" => DATA <= x"203c";
            when "01" & x"0e9" => DATA <= x"003f";
            when "01" & x"0ea" => DATA <= x"2b26";
            when "01" & x"0eb" => DATA <= x"6100";
            when "01" & x"0ec" => DATA <= x"e826";
            when "01" & x"0ed" => DATA <= x"6100";
            when "01" & x"0ee" => DATA <= x"e836";
            when "01" & x"0ef" => DATA <= x"21fc";
            when "01" & x"0f0" => DATA <= x"4430";
            when "01" & x"0f1" => DATA <= x"3a00";
            when "01" & x"0f2" => DATA <= x"0600";
            when "01" & x"0f3" => DATA <= x"223c";
            when "01" & x"0f4" => DATA <= x"0000";
            when "01" & x"0f5" => DATA <= x"0603";
            when "01" & x"0f6" => DATA <= x"243c";
            when "01" & x"0f7" => DATA <= x"0000";
            when "01" & x"0f8" => DATA <= x"00fc";
            when "01" & x"0f9" => DATA <= x"6100";
            when "01" & x"0fa" => DATA <= x"f4f2";
            when "01" & x"0fb" => DATA <= x"11fc";
            when "01" & x"0fc" => DATA <= x"0020";
            when "01" & x"0fd" => DATA <= x"060b";
            when "01" & x"0fe" => DATA <= x"21fc";
            when "01" & x"0ff" => DATA <= x"4431";
            when "01" & x"100" => DATA <= x"3a00";
            when "01" & x"101" => DATA <= x"060c";
            when "01" & x"102" => DATA <= x"2001";
            when "01" & x"103" => DATA <= x"223c";
            when "01" & x"104" => DATA <= x"0000";
            when "01" & x"105" => DATA <= x"060f";
            when "01" & x"106" => DATA <= x"243c";
            when "01" & x"107" => DATA <= x"0000";
            when "01" & x"108" => DATA <= x"00f4";
            when "01" & x"109" => DATA <= x"6100";
            when "01" & x"10a" => DATA <= x"f4d2";
            when "01" & x"10b" => DATA <= x"11fc";
            when "01" & x"10c" => DATA <= x"0020";
            when "01" & x"10d" => DATA <= x"0617";
            when "01" & x"10e" => DATA <= x"21fc";
            when "01" & x"10f" => DATA <= x"4432";
            when "01" & x"110" => DATA <= x"3a00";
            when "01" & x"111" => DATA <= x"0618";
            when "01" & x"112" => DATA <= x"2002";
            when "01" & x"113" => DATA <= x"223c";
            when "01" & x"114" => DATA <= x"0000";
            when "01" & x"115" => DATA <= x"061b";
            when "01" & x"116" => DATA <= x"243c";
            when "01" & x"117" => DATA <= x"0000";
            when "01" & x"118" => DATA <= x"00e8";
            when "01" & x"119" => DATA <= x"6100";
            when "01" & x"11a" => DATA <= x"f4b2";
            when "01" & x"11b" => DATA <= x"11fc";
            when "01" & x"11c" => DATA <= x"0020";
            when "01" & x"11d" => DATA <= x"0623";
            when "01" & x"11e" => DATA <= x"21fc";
            when "01" & x"11f" => DATA <= x"4433";
            when "01" & x"120" => DATA <= x"3a00";
            when "01" & x"121" => DATA <= x"0624";
            when "01" & x"122" => DATA <= x"2003";
            when "01" & x"123" => DATA <= x"223c";
            when "01" & x"124" => DATA <= x"0000";
            when "01" & x"125" => DATA <= x"0627";
            when "01" & x"126" => DATA <= x"243c";
            when "01" & x"127" => DATA <= x"0000";
            when "01" & x"128" => DATA <= x"00dc";
            when "01" & x"129" => DATA <= x"6100";
            when "01" & x"12a" => DATA <= x"f492";
            when "01" & x"12b" => DATA <= x"11fc";
            when "01" & x"12c" => DATA <= x"0020";
            when "01" & x"12d" => DATA <= x"062f";
            when "01" & x"12e" => DATA <= x"21fc";
            when "01" & x"12f" => DATA <= x"5352";
            when "01" & x"130" => DATA <= x"3a00";
            when "01" & x"131" => DATA <= x"0630";
            when "01" & x"132" => DATA <= x"223c";
            when "01" & x"133" => DATA <= x"0000";
            when "01" & x"134" => DATA <= x"0633";
            when "01" & x"135" => DATA <= x"243c";
            when "01" & x"136" => DATA <= x"0000";
            when "01" & x"137" => DATA <= x"00cd";
            when "01" & x"138" => DATA <= x"40c0";
            when "01" & x"139" => DATA <= x"6100";
            when "01" & x"13a" => DATA <= x"f6b4";
            when "01" & x"13b" => DATA <= x"11fc";
            when "01" & x"13c" => DATA <= x"0020";
            when "01" & x"13d" => DATA <= x"0643";
            when "01" & x"13e" => DATA <= x"21fc";
            when "01" & x"13f" => DATA <= x"2020";
            when "01" & x"140" => DATA <= x"0a0d";
            when "01" & x"141" => DATA <= x"0644";
            when "01" & x"142" => DATA <= x"21fc";
            when "01" & x"143" => DATA <= x"4434";
            when "01" & x"144" => DATA <= x"3a00";
            when "01" & x"145" => DATA <= x"0648";
            when "01" & x"146" => DATA <= x"2004";
            when "01" & x"147" => DATA <= x"223c";
            when "01" & x"148" => DATA <= x"0000";
            when "01" & x"149" => DATA <= x"064b";
            when "01" & x"14a" => DATA <= x"243c";
            when "01" & x"14b" => DATA <= x"0000";
            when "01" & x"14c" => DATA <= x"00b8";
            when "01" & x"14d" => DATA <= x"6100";
            when "01" & x"14e" => DATA <= x"f44a";
            when "01" & x"14f" => DATA <= x"11fc";
            when "01" & x"150" => DATA <= x"0020";
            when "01" & x"151" => DATA <= x"0653";
            when "01" & x"152" => DATA <= x"21fc";
            when "01" & x"153" => DATA <= x"4435";
            when "01" & x"154" => DATA <= x"3a00";
            when "01" & x"155" => DATA <= x"0654";
            when "01" & x"156" => DATA <= x"2005";
            when "01" & x"157" => DATA <= x"223c";
            when "01" & x"158" => DATA <= x"0000";
            when "01" & x"159" => DATA <= x"0657";
            when "01" & x"15a" => DATA <= x"243c";
            when "01" & x"15b" => DATA <= x"0000";
            when "01" & x"15c" => DATA <= x"00ac";
            when "01" & x"15d" => DATA <= x"6100";
            when "01" & x"15e" => DATA <= x"f42a";
            when "01" & x"15f" => DATA <= x"11fc";
            when "01" & x"160" => DATA <= x"0020";
            when "01" & x"161" => DATA <= x"065f";
            when "01" & x"162" => DATA <= x"21fc";
            when "01" & x"163" => DATA <= x"4436";
            when "01" & x"164" => DATA <= x"3a00";
            when "01" & x"165" => DATA <= x"0660";
            when "01" & x"166" => DATA <= x"2006";
            when "01" & x"167" => DATA <= x"223c";
            when "01" & x"168" => DATA <= x"0000";
            when "01" & x"169" => DATA <= x"0663";
            when "01" & x"16a" => DATA <= x"243c";
            when "01" & x"16b" => DATA <= x"0000";
            when "01" & x"16c" => DATA <= x"00a0";
            when "01" & x"16d" => DATA <= x"6100";
            when "01" & x"16e" => DATA <= x"f40a";
            when "01" & x"16f" => DATA <= x"11fc";
            when "01" & x"170" => DATA <= x"0020";
            when "01" & x"171" => DATA <= x"066b";
            when "01" & x"172" => DATA <= x"21fc";
            when "01" & x"173" => DATA <= x"4437";
            when "01" & x"174" => DATA <= x"3a00";
            when "01" & x"175" => DATA <= x"066c";
            when "01" & x"176" => DATA <= x"2007";
            when "01" & x"177" => DATA <= x"223c";
            when "01" & x"178" => DATA <= x"0000";
            when "01" & x"179" => DATA <= x"066f";
            when "01" & x"17a" => DATA <= x"243c";
            when "01" & x"17b" => DATA <= x"0000";
            when "01" & x"17c" => DATA <= x"0094";
            when "01" & x"17d" => DATA <= x"6100";
            when "01" & x"17e" => DATA <= x"f3ea";
            when "01" & x"17f" => DATA <= x"11fc";
            when "01" & x"180" => DATA <= x"0020";
            when "01" & x"181" => DATA <= x"0677";
            when "01" & x"182" => DATA <= x"21fc";
            when "01" & x"183" => DATA <= x"5553";
            when "01" & x"184" => DATA <= x"3a00";
            when "01" & x"185" => DATA <= x"0678";
            when "01" & x"186" => DATA <= x"4e68";
            when "01" & x"187" => DATA <= x"2008";
            when "01" & x"188" => DATA <= x"223c";
            when "01" & x"189" => DATA <= x"0000";
            when "01" & x"18a" => DATA <= x"067b";
            when "01" & x"18b" => DATA <= x"243c";
            when "01" & x"18c" => DATA <= x"0000";
            when "01" & x"18d" => DATA <= x"0094";
            when "01" & x"18e" => DATA <= x"6100";
            when "01" & x"18f" => DATA <= x"f3c8";
            when "01" & x"190" => DATA <= x"11fc";
            when "01" & x"191" => DATA <= x"0020";
            when "01" & x"192" => DATA <= x"0683";
            when "01" & x"193" => DATA <= x"21fc";
            when "01" & x"194" => DATA <= x"2020";
            when "01" & x"195" => DATA <= x"0a0d";
            when "01" & x"196" => DATA <= x"0684";
            when "01" & x"197" => DATA <= x"21fc";
            when "01" & x"198" => DATA <= x"4130";
            when "01" & x"199" => DATA <= x"3a00";
            when "01" & x"19a" => DATA <= x"0688";
            when "01" & x"19b" => DATA <= x"2008";
            when "01" & x"19c" => DATA <= x"223c";
            when "01" & x"19d" => DATA <= x"0000";
            when "01" & x"19e" => DATA <= x"068b";
            when "01" & x"19f" => DATA <= x"243c";
            when "01" & x"1a0" => DATA <= x"0000";
            when "01" & x"1a1" => DATA <= x"0094";
            when "01" & x"1a2" => DATA <= x"6100";
            when "01" & x"1a3" => DATA <= x"f3a0";
            when "01" & x"1a4" => DATA <= x"11fc";
            when "01" & x"1a5" => DATA <= x"0020";
            when "01" & x"1a6" => DATA <= x"0693";
            when "01" & x"1a7" => DATA <= x"21fc";
            when "01" & x"1a8" => DATA <= x"4131";
            when "01" & x"1a9" => DATA <= x"3a00";
            when "01" & x"1aa" => DATA <= x"0694";
            when "01" & x"1ab" => DATA <= x"2009";
            when "01" & x"1ac" => DATA <= x"223c";
            when "01" & x"1ad" => DATA <= x"0000";
            when "01" & x"1ae" => DATA <= x"0697";
            when "01" & x"1af" => DATA <= x"243c";
            when "01" & x"1b0" => DATA <= x"0000";
            when "01" & x"1b1" => DATA <= x"0094";
            when "01" & x"1b2" => DATA <= x"6100";
            when "01" & x"1b3" => DATA <= x"f380";
            when "01" & x"1b4" => DATA <= x"11fc";
            when "01" & x"1b5" => DATA <= x"0020";
            when "01" & x"1b6" => DATA <= x"069f";
            when "01" & x"1b7" => DATA <= x"21fc";
            when "01" & x"1b8" => DATA <= x"4132";
            when "01" & x"1b9" => DATA <= x"3a00";
            when "01" & x"1ba" => DATA <= x"06a0";
            when "01" & x"1bb" => DATA <= x"200a";
            when "01" & x"1bc" => DATA <= x"223c";
            when "01" & x"1bd" => DATA <= x"0000";
            when "01" & x"1be" => DATA <= x"06a3";
            when "01" & x"1bf" => DATA <= x"243c";
            when "01" & x"1c0" => DATA <= x"0000";
            when "01" & x"1c1" => DATA <= x"0094";
            when "01" & x"1c2" => DATA <= x"6100";
            when "01" & x"1c3" => DATA <= x"f360";
            when "01" & x"1c4" => DATA <= x"11fc";
            when "01" & x"1c5" => DATA <= x"0020";
            when "01" & x"1c6" => DATA <= x"06ab";
            when "01" & x"1c7" => DATA <= x"21fc";
            when "01" & x"1c8" => DATA <= x"4133";
            when "01" & x"1c9" => DATA <= x"3a00";
            when "01" & x"1ca" => DATA <= x"06ac";
            when "01" & x"1cb" => DATA <= x"200b";
            when "01" & x"1cc" => DATA <= x"223c";
            when "01" & x"1cd" => DATA <= x"0000";
            when "01" & x"1ce" => DATA <= x"06af";
            when "01" & x"1cf" => DATA <= x"243c";
            when "01" & x"1d0" => DATA <= x"0000";
            when "01" & x"1d1" => DATA <= x"0094";
            when "01" & x"1d2" => DATA <= x"6100";
            when "01" & x"1d3" => DATA <= x"f340";
            when "01" & x"1d4" => DATA <= x"11fc";
            when "01" & x"1d5" => DATA <= x"0020";
            when "01" & x"1d6" => DATA <= x"06b7";
            when "01" & x"1d7" => DATA <= x"21fc";
            when "01" & x"1d8" => DATA <= x"5353";
            when "01" & x"1d9" => DATA <= x"3a00";
            when "01" & x"1da" => DATA <= x"06b8";
            when "01" & x"1db" => DATA <= x"200f";
            when "01" & x"1dc" => DATA <= x"223c";
            when "01" & x"1dd" => DATA <= x"0000";
            when "01" & x"1de" => DATA <= x"06bb";
            when "01" & x"1df" => DATA <= x"243c";
            when "01" & x"1e0" => DATA <= x"0000";
            when "01" & x"1e1" => DATA <= x"0094";
            when "01" & x"1e2" => DATA <= x"6100";
            when "01" & x"1e3" => DATA <= x"f320";
            when "01" & x"1e4" => DATA <= x"11fc";
            when "01" & x"1e5" => DATA <= x"0020";
            when "01" & x"1e6" => DATA <= x"06c3";
            when "01" & x"1e7" => DATA <= x"21fc";
            when "01" & x"1e8" => DATA <= x"2020";
            when "01" & x"1e9" => DATA <= x"0a0d";
            when "01" & x"1ea" => DATA <= x"06c4";
            when "01" & x"1eb" => DATA <= x"21fc";
            when "01" & x"1ec" => DATA <= x"4134";
            when "01" & x"1ed" => DATA <= x"3a00";
            when "01" & x"1ee" => DATA <= x"06c8";
            when "01" & x"1ef" => DATA <= x"200c";
            when "01" & x"1f0" => DATA <= x"223c";
            when "01" & x"1f1" => DATA <= x"0000";
            when "01" & x"1f2" => DATA <= x"06cb";
            when "01" & x"1f3" => DATA <= x"243c";
            when "01" & x"1f4" => DATA <= x"0000";
            when "01" & x"1f5" => DATA <= x"0094";
            when "01" & x"1f6" => DATA <= x"6100";
            when "01" & x"1f7" => DATA <= x"f2f8";
            when "01" & x"1f8" => DATA <= x"11fc";
            when "01" & x"1f9" => DATA <= x"0020";
            when "01" & x"1fa" => DATA <= x"06d3";
            when "01" & x"1fb" => DATA <= x"21fc";
            when "01" & x"1fc" => DATA <= x"4135";
            when "01" & x"1fd" => DATA <= x"3a00";
            when "01" & x"1fe" => DATA <= x"06d4";
            when "01" & x"1ff" => DATA <= x"200d";
            when "01" & x"200" => DATA <= x"223c";
            when "01" & x"201" => DATA <= x"0000";
            when "01" & x"202" => DATA <= x"06d7";
            when "01" & x"203" => DATA <= x"243c";
            when "01" & x"204" => DATA <= x"0000";
            when "01" & x"205" => DATA <= x"0094";
            when "01" & x"206" => DATA <= x"6100";
            when "01" & x"207" => DATA <= x"f2d8";
            when "01" & x"208" => DATA <= x"11fc";
            when "01" & x"209" => DATA <= x"0020";
            when "01" & x"20a" => DATA <= x"06df";
            when "01" & x"20b" => DATA <= x"21fc";
            when "01" & x"20c" => DATA <= x"4136";
            when "01" & x"20d" => DATA <= x"3a00";
            when "01" & x"20e" => DATA <= x"06e0";
            when "01" & x"20f" => DATA <= x"200e";
            when "01" & x"210" => DATA <= x"223c";
            when "01" & x"211" => DATA <= x"0000";
            when "01" & x"212" => DATA <= x"06e3";
            when "01" & x"213" => DATA <= x"243c";
            when "01" & x"214" => DATA <= x"0000";
            when "01" & x"215" => DATA <= x"0094";
            when "01" & x"216" => DATA <= x"6100";
            when "01" & x"217" => DATA <= x"f2b8";
            when "01" & x"218" => DATA <= x"11fc";
            when "01" & x"219" => DATA <= x"0020";
            when "01" & x"21a" => DATA <= x"06eb";
            when "01" & x"21b" => DATA <= x"21fc";
            when "01" & x"21c" => DATA <= x"4137";
            when "01" & x"21d" => DATA <= x"3a00";
            when "01" & x"21e" => DATA <= x"06ec";
            when "01" & x"21f" => DATA <= x"200f";
            when "01" & x"220" => DATA <= x"223c";
            when "01" & x"221" => DATA <= x"0000";
            when "01" & x"222" => DATA <= x"06ef";
            when "01" & x"223" => DATA <= x"243c";
            when "01" & x"224" => DATA <= x"0000";
            when "01" & x"225" => DATA <= x"0094";
            when "01" & x"226" => DATA <= x"6100";
            when "01" & x"227" => DATA <= x"f298";
            when "01" & x"228" => DATA <= x"11fc";
            when "01" & x"229" => DATA <= x"0020";
            when "01" & x"22a" => DATA <= x"06f7";
            when "01" & x"22b" => DATA <= x"21fc";
            when "01" & x"22c" => DATA <= x"5043";
            when "01" & x"22d" => DATA <= x"3a00";
            when "01" & x"22e" => DATA <= x"06f8";
            when "01" & x"22f" => DATA <= x"203c";
            when "01" & x"230" => DATA <= x"0000";
            when "01" & x"231" => DATA <= x"0600";
            when "01" & x"232" => DATA <= x"6100";
            when "01" & x"233" => DATA <= x"e598";
            when "01" & x"234" => DATA <= x"6100";
            when "01" & x"235" => DATA <= x"e5a8";
            when "01" & x"236" => DATA <= x"6000";
            when "01" & x"237" => DATA <= x"f956";
            when "01" & x"238" => DATA <= x"203c";
            when "01" & x"239" => DATA <= x"003f";
            when "01" & x"23a" => DATA <= x"2945";
            when "01" & x"23b" => DATA <= x"6100";
            when "01" & x"23c" => DATA <= x"e586";
            when "01" & x"23d" => DATA <= x"4e75";
            when "01" & x"23e" => DATA <= x"6000";
            when "01" & x"23f" => DATA <= x"e9c6";
            when "01" & x"240" => DATA <= x"6000";
            when "01" & x"241" => DATA <= x"e2f4";
            when "01" & x"242" => DATA <= x"7010";
            when "01" & x"243" => DATA <= x"220e";
            when "01" & x"244" => DATA <= x"6100";
            when "01" & x"245" => DATA <= x"eb42";
            when "01" & x"246" => DATA <= x"6900";
            when "01" & x"247" => DATA <= x"00d2";
            when "01" & x"248" => DATA <= x"2e02";
            when "01" & x"249" => DATA <= x"6100";
            when "01" & x"24a" => DATA <= x"029a";
            when "01" & x"24b" => DATA <= x"7010";
            when "01" & x"24c" => DATA <= x"6100";
            when "01" & x"24d" => DATA <= x"eb32";
            when "01" & x"24e" => DATA <= x"6900";
            when "01" & x"24f" => DATA <= x"00c2";
            when "01" & x"250" => DATA <= x"2c02";
            when "01" & x"251" => DATA <= x"6100";
            when "01" & x"252" => DATA <= x"028a";
            when "01" & x"253" => DATA <= x"7010";
            when "01" & x"254" => DATA <= x"6100";
            when "01" & x"255" => DATA <= x"eb22";
            when "01" & x"256" => DATA <= x"6900";
            when "01" & x"257" => DATA <= x"00b2";
            when "01" & x"258" => DATA <= x"2c41";
            when "01" & x"259" => DATA <= x"2a02";
            when "01" & x"25a" => DATA <= x"6100";
            when "01" & x"25b" => DATA <= x"026a";
            when "01" & x"25c" => DATA <= x"101e";
            when "01" & x"25d" => DATA <= x"0200";
            when "01" & x"25e" => DATA <= x"00df";
            when "01" & x"25f" => DATA <= x"b03c";
            when "01" & x"260" => DATA <= x"0052";
            when "01" & x"261" => DATA <= x"6700";
            when "01" & x"262" => DATA <= x"0012";
            when "01" & x"263" => DATA <= x"b03c";
            when "01" & x"264" => DATA <= x"0057";
            when "01" & x"265" => DATA <= x"6600";
            when "01" & x"266" => DATA <= x"0094";
            when "01" & x"267" => DATA <= x"183c";
            when "01" & x"268" => DATA <= x"0006";
            when "01" & x"269" => DATA <= x"6000";
            when "01" & x"26a" => DATA <= x"0006";
            when "01" & x"26b" => DATA <= x"183c";
            when "01" & x"26c" => DATA <= x"0007";
            when "01" & x"26d" => DATA <= x"6100";
            when "01" & x"26e" => DATA <= x"0244";
            when "01" & x"26f" => DATA <= x"6700";
            when "01" & x"270" => DATA <= x"0020";
            when "01" & x"271" => DATA <= x"101e";
            when "01" & x"272" => DATA <= x"0200";
            when "01" & x"273" => DATA <= x"00df";
            when "01" & x"274" => DATA <= x"b03c";
            when "01" & x"275" => DATA <= x"0053";
            when "01" & x"276" => DATA <= x"6700";
            when "01" & x"277" => DATA <= x"001a";
            when "01" & x"278" => DATA <= x"b03c";
            when "01" & x"279" => DATA <= x"004d";
            when "01" & x"27a" => DATA <= x"6600";
            when "01" & x"27b" => DATA <= x"006a";
            when "01" & x"27c" => DATA <= x"163c";
            when "01" & x"27d" => DATA <= x"0040";
            when "01" & x"27e" => DATA <= x"6000";
            when "01" & x"27f" => DATA <= x"000e";
            when "01" & x"280" => DATA <= x"103c";
            when "01" & x"281" => DATA <= x"0010";
            when "01" & x"282" => DATA <= x"6000";
            when "01" & x"283" => DATA <= x"0006";
            when "01" & x"284" => DATA <= x"163c";
            when "01" & x"285" => DATA <= x"0020";
            when "01" & x"286" => DATA <= x"6100";
            when "01" & x"287" => DATA <= x"0212";
            when "01" & x"288" => DATA <= x"6600";
            when "01" & x"289" => DATA <= x"f798";
            when "01" & x"28a" => DATA <= x"11fc";
            when "01" & x"28b" => DATA <= x"000e";
            when "01" & x"28c" => DATA <= x"0600";
            when "01" & x"28d" => DATA <= x"11fc";
            when "01" & x"28e" => DATA <= x"0010";
            when "01" & x"28f" => DATA <= x"0601";
            when "01" & x"290" => DATA <= x"21c7";
            when "01" & x"291" => DATA <= x"0602";
            when "01" & x"292" => DATA <= x"21c6";
            when "01" & x"293" => DATA <= x"0606";
            when "01" & x"294" => DATA <= x"31c5";
            when "01" & x"295" => DATA <= x"060a";
            when "01" & x"296" => DATA <= x"11c4";
            when "01" & x"297" => DATA <= x"060c";
            when "01" & x"298" => DATA <= x"11c3";
            when "01" & x"299" => DATA <= x"060d";
            when "01" & x"29a" => DATA <= x"223c";
            when "01" & x"29b" => DATA <= x"0000";
            when "01" & x"29c" => DATA <= x"0600";
            when "01" & x"29d" => DATA <= x"203c";
            when "01" & x"29e" => DATA <= x"0000";
            when "01" & x"29f" => DATA <= x"00fa";
            when "01" & x"2a0" => DATA <= x"6100";
            when "01" & x"2a1" => DATA <= x"e6a2";
            when "01" & x"2a2" => DATA <= x"0c04";
            when "01" & x"2a3" => DATA <= x"0006";
            when "01" & x"2a4" => DATA <= x"6600";
            when "01" & x"2a5" => DATA <= x"000c";
            when "01" & x"2a6" => DATA <= x"2a47";
            when "01" & x"2a7" => DATA <= x"2c46";
            when "01" & x"2a8" => DATA <= x"2405";
            when "01" & x"2a9" => DATA <= x"6000";
            when "01" & x"2aa" => DATA <= x"014c";
            when "01" & x"2ab" => DATA <= x"2a46";
            when "01" & x"2ac" => DATA <= x"2c47";
            when "01" & x"2ad" => DATA <= x"2405";
            when "01" & x"2ae" => DATA <= x"6000";
            when "01" & x"2af" => DATA <= x"015c";
            when "01" & x"2b0" => DATA <= x"203c";
            when "01" & x"2b1" => DATA <= x"003f";
            when "01" & x"2b2" => DATA <= x"2969";
            when "01" & x"2b3" => DATA <= x"6100";
            when "01" & x"2b4" => DATA <= x"e496";
            when "01" & x"2b5" => DATA <= x"4e75";
            when "01" & x"2b6" => DATA <= x"6100";
            when "01" & x"2b7" => DATA <= x"e4a4";
            when "01" & x"2b8" => DATA <= x"5880";
            when "01" & x"2b9" => DATA <= x"6100";
            when "01" & x"2ba" => DATA <= x"e48a";
            when "01" & x"2bb" => DATA <= x"0cb8";
            when "01" & x"2bc" => DATA <= x"0000";
            when "01" & x"2bd" => DATA <= x"0000";
            when "01" & x"2be" => DATA <= x"0510";
            when "01" & x"2bf" => DATA <= x"6700";
            when "01" & x"2c0" => DATA <= x"0022";
            when "01" & x"2c1" => DATA <= x"203c";
            when "01" & x"2c2" => DATA <= x"003f";
            when "01" & x"2c3" => DATA <= x"2c54";
            when "01" & x"2c4" => DATA <= x"6100";
            when "01" & x"2c5" => DATA <= x"e474";
            when "01" & x"2c6" => DATA <= x"2038";
            when "01" & x"2c7" => DATA <= x"0510";
            when "01" & x"2c8" => DATA <= x"223c";
            when "01" & x"2c9" => DATA <= x"0000";
            when "01" & x"2ca" => DATA <= x"0600";
            when "01" & x"2cb" => DATA <= x"143c";
            when "01" & x"2cc" => DATA <= x"00ff";
            when "01" & x"2cd" => DATA <= x"6100";
            when "01" & x"2ce" => DATA <= x"f14a";
            when "01" & x"2cf" => DATA <= x"6100";
            when "01" & x"2d0" => DATA <= x"e45e";
            when "01" & x"2d1" => DATA <= x"6100";
            when "01" & x"2d2" => DATA <= x"e46e";
            when "01" & x"2d3" => DATA <= x"2e78";
            when "01" & x"2d4" => DATA <= x"0508";
            when "01" & x"2d5" => DATA <= x"6000";
            when "01" & x"2d6" => DATA <= x"ddb2";
            when "01" & x"2d7" => DATA <= x"2f00";
            when "01" & x"2d8" => DATA <= x"203c";
            when "01" & x"2d9" => DATA <= x"003f";
            when "01" & x"2da" => DATA <= x"2d18";
            when "01" & x"2db" => DATA <= x"21fc";
            when "01" & x"2dc" => DATA <= x"0000";
            when "01" & x"2dd" => DATA <= x"0000";
            when "01" & x"2de" => DATA <= x"0510";
            when "01" & x"2df" => DATA <= x"6100";
            when "01" & x"2e0" => DATA <= x"eb60";
            when "01" & x"2e1" => DATA <= x"201f";
            when "01" & x"2e2" => DATA <= x"4e75";
            when "01" & x"2e3" => DATA <= x"0839";
            when "01" & x"2e4" => DATA <= x"0006";
            when "01" & x"2e5" => DATA <= x"fffe";
            when "01" & x"2e6" => DATA <= x"0000";
            when "01" & x"2e7" => DATA <= x"67f6";
            when "01" & x"2e8" => DATA <= x"13c0";
            when "01" & x"2e9" => DATA <= x"fffe";
            when "01" & x"2ea" => DATA <= x"0001";
            when "01" & x"2eb" => DATA <= x"4e75";
            when "01" & x"2ec" => DATA <= x"4e75";
            when "01" & x"2ed" => DATA <= x"2f00";
            when "01" & x"2ee" => DATA <= x"203c";
            when "01" & x"2ef" => DATA <= x"003f";
            when "01" & x"2f0" => DATA <= x"2e38";
            when "01" & x"2f1" => DATA <= x"6100";
            when "01" & x"2f2" => DATA <= x"eb3c";
            when "01" & x"2f3" => DATA <= x"201f";
            when "01" & x"2f4" => DATA <= x"4e75";
            when "01" & x"2f5" => DATA <= x"b07c";
            when "01" & x"2f6" => DATA <= x"0010";
            when "01" & x"2f7" => DATA <= x"6300";
            when "01" & x"2f8" => DATA <= x"000e";
            when "01" & x"2f9" => DATA <= x"203c";
            when "01" & x"2fa" => DATA <= x"003f";
            when "01" & x"2fb" => DATA <= x"2e1c";
            when "01" & x"2fc" => DATA <= x"003c";
            when "01" & x"2fd" => DATA <= x"0002";
            when "01" & x"2fe" => DATA <= x"4e75";
            when "01" & x"2ff" => DATA <= x"41f9";
            when "01" & x"300" => DATA <= x"003f";
            when "01" & x"301" => DATA <= x"362c";
            when "01" & x"302" => DATA <= x"e588";
            when "01" & x"303" => DATA <= x"d1c0";
            when "01" & x"304" => DATA <= x"d1c0";
            when "01" & x"305" => DATA <= x"d1c0";
            when "01" & x"306" => DATA <= x"2258";
            when "01" & x"307" => DATA <= x"b3fc";
            when "01" & x"308" => DATA <= x"0000";
            when "01" & x"309" => DATA <= x"0000";
            when "01" & x"30a" => DATA <= x"67dc";
            when "01" & x"30b" => DATA <= x"2f04";
            when "01" & x"30c" => DATA <= x"2458";
            when "01" & x"30d" => DATA <= x"2658";
            when "01" & x"30e" => DATA <= x"4a81";
            when "01" & x"30f" => DATA <= x"6600";
            when "01" & x"310" => DATA <= x"0008";
            when "01" & x"311" => DATA <= x"2211";
            when "01" & x"312" => DATA <= x"6000";
            when "01" & x"313" => DATA <= x"0008";
            when "01" & x"314" => DATA <= x"2811";
            when "01" & x"315" => DATA <= x"2281";
            when "01" & x"316" => DATA <= x"c941";
            when "01" & x"317" => DATA <= x"4a82";
            when "01" & x"318" => DATA <= x"6600";
            when "01" & x"319" => DATA <= x"0008";
            when "01" & x"31a" => DATA <= x"2412";
            when "01" & x"31b" => DATA <= x"6000";
            when "01" & x"31c" => DATA <= x"0008";
            when "01" & x"31d" => DATA <= x"2812";
            when "01" & x"31e" => DATA <= x"2482";
            when "01" & x"31f" => DATA <= x"c942";
            when "01" & x"320" => DATA <= x"4a83";
            when "01" & x"321" => DATA <= x"6600";
            when "01" & x"322" => DATA <= x"0008";
            when "01" & x"323" => DATA <= x"2612";
            when "01" & x"324" => DATA <= x"6000";
            when "01" & x"325" => DATA <= x"0008";
            when "01" & x"326" => DATA <= x"2813";
            when "01" & x"327" => DATA <= x"2681";
            when "01" & x"328" => DATA <= x"c941";
            when "01" & x"329" => DATA <= x"281f";
            when "01" & x"32a" => DATA <= x"4e75";
            when "01" & x"32b" => DATA <= x"6000";
            when "01" & x"32c" => DATA <= x"e11e";
            when "01" & x"32d" => DATA <= x"6000";
            when "01" & x"32e" => DATA <= x"e11a";
            when "01" & x"32f" => DATA <= x"0200";
            when "01" & x"330" => DATA <= x"0040";
            when "01" & x"331" => DATA <= x"8138";
            when "01" & x"332" => DATA <= x"0535";
            when "01" & x"333" => DATA <= x"4e75";
            when "01" & x"334" => DATA <= x"21fc";
            when "01" & x"335" => DATA <= x"0000";
            when "01" & x"336" => DATA <= x"0000";
            when "01" & x"337" => DATA <= x"0518";
            when "01" & x"338" => DATA <= x"b2bc";
            when "01" & x"339" => DATA <= x"4142";
            when "01" & x"33a" => DATA <= x"4558";
            when "01" & x"33b" => DATA <= x"6600";
            when "01" & x"33c" => DATA <= x"0018";
            when "01" & x"33d" => DATA <= x"21c2";
            when "01" & x"33e" => DATA <= x"0518";
            when "01" & x"33f" => DATA <= x"b4b8";
            when "01" & x"340" => DATA <= x"051c";
            when "01" & x"341" => DATA <= x"6300";
            when "01" & x"342" => DATA <= x"000c";
            when "01" & x"343" => DATA <= x"203c";
            when "01" & x"344" => DATA <= x"003f";
            when "01" & x"345" => DATA <= x"2e60";
            when "01" & x"346" => DATA <= x"6100";
            when "01" & x"347" => DATA <= x"ea92";
            when "01" & x"348" => DATA <= x"2e78";
            when "01" & x"349" => DATA <= x"0508";
            when "01" & x"34a" => DATA <= x"6000";
            when "01" & x"34b" => DATA <= x"dcc8";
            when "01" & x"34c" => DATA <= x"6000";
            when "01" & x"34d" => DATA <= x"e0dc";
            when "01" & x"34e" => DATA <= x"6000";
            when "01" & x"34f" => DATA <= x"e0d8";
            when "01" & x"350" => DATA <= x"21cd";
            when "01" & x"351" => DATA <= x"0600";
            when "01" & x"352" => DATA <= x"223c";
            when "01" & x"353" => DATA <= x"0000";
            when "01" & x"354" => DATA <= x"0600";
            when "01" & x"355" => DATA <= x"7005";
            when "01" & x"356" => DATA <= x"6100";
            when "01" & x"357" => DATA <= x"e536";
            when "01" & x"358" => DATA <= x"1cf8";
            when "01" & x"359" => DATA <= x"0605";
            when "01" & x"35a" => DATA <= x"51ca";
            when "01" & x"35b" => DATA <= x"ffee";
            when "01" & x"35c" => DATA <= x"4e75";
            when "01" & x"35d" => DATA <= x"21cd";
            when "01" & x"35e" => DATA <= x"0600";
            when "01" & x"35f" => DATA <= x"223c";
            when "01" & x"360" => DATA <= x"0000";
            when "01" & x"361" => DATA <= x"0600";
            when "01" & x"362" => DATA <= x"11de";
            when "01" & x"363" => DATA <= x"0605";
            when "01" & x"364" => DATA <= x"7006";
            when "01" & x"365" => DATA <= x"6100";
            when "01" & x"366" => DATA <= x"e518";
            when "01" & x"367" => DATA <= x"51ca";
            when "01" & x"368" => DATA <= x"ffee";
            when "01" & x"369" => DATA <= x"4e75";
            when "01" & x"36a" => DATA <= x"2a7c";
            when "01" & x"36b" => DATA <= x"003f";
            when "01" & x"36c" => DATA <= x"37e4";
            when "01" & x"36d" => DATA <= x"2c7c";
            when "01" & x"36e" => DATA <= x"ffff";
            when "01" & x"36f" => DATA <= x"2500";
            when "01" & x"370" => DATA <= x"243c";
            when "01" & x"371" => DATA <= x"0000";
            when "01" & x"372" => DATA <= x"01fb";
            when "01" & x"373" => DATA <= x"61d2";
            when "01" & x"374" => DATA <= x"2a7c";
            when "01" & x"375" => DATA <= x"ffff";
            when "01" & x"376" => DATA <= x"0200";
            when "01" & x"377" => DATA <= x"2c7c";
            when "01" & x"378" => DATA <= x"0000";
            when "01" & x"379" => DATA <= x"0600";
            when "01" & x"37a" => DATA <= x"7402";
            when "01" & x"37b" => DATA <= x"61a8";
            when "01" & x"37c" => DATA <= x"2a7c";
            when "01" & x"37d" => DATA <= x"0000";
            when "01" & x"37e" => DATA <= x"0600";
            when "01" & x"37f" => DATA <= x"2c7c";
            when "01" & x"380" => DATA <= x"ffff";
            when "01" & x"381" => DATA <= x"2503";
            when "01" & x"382" => DATA <= x"7402";
            when "01" & x"383" => DATA <= x"61b2";
            when "01" & x"384" => DATA <= x"31fc";
            when "01" & x"385" => DATA <= x"2500";
            when "01" & x"386" => DATA <= x"0600";
            when "01" & x"387" => DATA <= x"2a7c";
            when "01" & x"388" => DATA <= x"0000";
            when "01" & x"389" => DATA <= x"0600";
            when "01" & x"38a" => DATA <= x"2c7c";
            when "01" & x"38b" => DATA <= x"ffff";
            when "01" & x"38c" => DATA <= x"0200";
            when "01" & x"38d" => DATA <= x"7402";
            when "01" & x"38e" => DATA <= x"619c";
            when "01" & x"38f" => DATA <= x"4e75";
            when "01" & x"390" => DATA <= x"0c1e";
            when "01" & x"391" => DATA <= x"0020";
            when "01" & x"392" => DATA <= x"67fa";
            when "01" & x"393" => DATA <= x"1026";
            when "01" & x"394" => DATA <= x"b03c";
            when "01" & x"395" => DATA <= x"000d";
            when "01" & x"396" => DATA <= x"4e75";
            when "01" & x"397" => DATA <= x"c38e";
            when "01" & x"398" => DATA <= x"0c1e";
            when "01" & x"399" => DATA <= x"0020";
            when "01" & x"39a" => DATA <= x"67fa";
            when "01" & x"39b" => DATA <= x"1026";
            when "01" & x"39c" => DATA <= x"c38e";
            when "01" & x"39d" => DATA <= x"b03c";
            when "01" & x"39e" => DATA <= x"000d";
            when "01" & x"39f" => DATA <= x"4e75";
            when "01" & x"3a0" => DATA <= x"7010";
            when "01" & x"3a1" => DATA <= x"220e";
            when "01" & x"3a2" => DATA <= x"6100";
            when "01" & x"3a3" => DATA <= x"e886";
            when "01" & x"3a4" => DATA <= x"6900";
            when "01" & x"3a5" => DATA <= x"000c";
            when "01" & x"3a6" => DATA <= x"2c41";
            when "01" & x"3a7" => DATA <= x"2202";
            when "01" & x"3a8" => DATA <= x"023c";
            when "01" & x"3a9" => DATA <= x"00fe";
            when "01" & x"3aa" => DATA <= x"4e75";
            when "01" & x"3ab" => DATA <= x"2c41";
            when "01" & x"3ac" => DATA <= x"2202";
            when "01" & x"3ad" => DATA <= x"003c";
            when "01" & x"3ae" => DATA <= x"0001";
            when "01" & x"3af" => DATA <= x"4e75";
            when "01" & x"3b0" => DATA <= x"4281";
            when "01" & x"3b1" => DATA <= x"101e";
            when "01" & x"3b2" => DATA <= x"2f00";
            when "01" & x"3b3" => DATA <= x"0c00";
            when "01" & x"3b4" => DATA <= x"0030";
            when "01" & x"3b5" => DATA <= x"6500";
            when "01" & x"3b6" => DATA <= x"002c";
            when "01" & x"3b7" => DATA <= x"0c00";
            when "01" & x"3b8" => DATA <= x"0039";
            when "01" & x"3b9" => DATA <= x"6300";
            when "01" & x"3ba" => DATA <= x"0018";
            when "01" & x"3bb" => DATA <= x"0200";
            when "01" & x"3bc" => DATA <= x"00df";
            when "01" & x"3bd" => DATA <= x"0c00";
            when "01" & x"3be" => DATA <= x"0041";
            when "01" & x"3bf" => DATA <= x"6500";
            when "01" & x"3c0" => DATA <= x"0018";
            when "01" & x"3c1" => DATA <= x"0c00";
            when "01" & x"3c2" => DATA <= x"0046";
            when "01" & x"3c3" => DATA <= x"6200";
            when "01" & x"3c4" => DATA <= x"0010";
            when "01" & x"3c5" => DATA <= x"5f00";
            when "01" & x"3c6" => DATA <= x"0200";
            when "01" & x"3c7" => DATA <= x"000f";
            when "01" & x"3c8" => DATA <= x"e981";
            when "01" & x"3c9" => DATA <= x"d200";
            when "01" & x"3ca" => DATA <= x"201f";
            when "01" & x"3cb" => DATA <= x"60ca";
            when "01" & x"3cc" => DATA <= x"201f";
            when "01" & x"3cd" => DATA <= x"0c00";
            when "01" & x"3ce" => DATA <= x"000d";
            when "01" & x"3cf" => DATA <= x"6700";
            when "01" & x"3d0" => DATA <= x"0012";
            when "01" & x"3d1" => DATA <= x"0c00";
            when "01" & x"3d2" => DATA <= x"0020";
            when "01" & x"3d3" => DATA <= x"6700";
            when "01" & x"3d4" => DATA <= x"000a";
            when "01" & x"3d5" => DATA <= x"534e";
            when "01" & x"3d6" => DATA <= x"003c";
            when "01" & x"3d7" => DATA <= x"0001";
            when "01" & x"3d8" => DATA <= x"4e75";
            when "01" & x"3d9" => DATA <= x"534e";
            when "01" & x"3da" => DATA <= x"023c";
            when "01" & x"3db" => DATA <= x"00fe";
            when "01" & x"3dc" => DATA <= x"4e75";
            when "01" & x"3dd" => DATA <= x"101e";
            when "01" & x"3de" => DATA <= x"0c00";
            when "01" & x"3df" => DATA <= x"0020";
            when "01" & x"3e0" => DATA <= x"6500";
            when "01" & x"3e1" => DATA <= x"000a";
            when "01" & x"3e2" => DATA <= x"0c00";
            when "01" & x"3e3" => DATA <= x"007f";
            when "01" & x"3e4" => DATA <= x"6500";
            when "01" & x"3e5" => DATA <= x"0006";
            when "01" & x"3e6" => DATA <= x"103c";
            when "01" & x"3e7" => DATA <= x"002e";
            when "01" & x"3e8" => DATA <= x"4e75";
            when "01" & x"3e9" => DATA <= x"0280";
            when "01" & x"3ea" => DATA <= x"0000";
            when "01" & x"3eb" => DATA <= x"0007";
            when "01" & x"3ec" => DATA <= x"e140";
            when "01" & x"3ed" => DATA <= x"027c";
            when "01" & x"3ee" => DATA <= x"f8ff";
            when "01" & x"3ef" => DATA <= x"221f";
            when "01" & x"3f0" => DATA <= x"4e75";
            when "01" & x"3f1" => DATA <= x"0d0a";
            when "01" & x"3f2" => DATA <= x"4163";
            when "01" & x"3f3" => DATA <= x"6f72";
            when "01" & x"3f4" => DATA <= x"6e20";
            when "01" & x"3f5" => DATA <= x"3638";
            when "01" & x"3f6" => DATA <= x"0020";
            when "01" & x"3f7" => DATA <= x"7365";
            when "01" & x"3f8" => DATA <= x"636f";
            when "01" & x"3f9" => DATA <= x"6e64";
            when "01" & x"3fa" => DATA <= x"2070";
            when "01" & x"3fb" => DATA <= x"726f";
            when "01" & x"3fc" => DATA <= x"6365";
            when "01" & x"3fd" => DATA <= x"7373";
            when "01" & x"3fe" => DATA <= x"6f72";
            when "01" & x"3ff" => DATA <= x"2000";
            when "01" & x"400" => DATA <= x"3030";
            when "01" & x"401" => DATA <= x"3830";
            when "01" & x"402" => DATA <= x"3030";
            when "01" & x"403" => DATA <= x"3031";
            when "01" & x"404" => DATA <= x"3030";
            when "01" & x"405" => DATA <= x"3230";
            when "01" & x"406" => DATA <= x"3033";
            when "01" & x"407" => DATA <= x"3030";
            when "01" & x"408" => DATA <= x"3430";
            when "01" & x"409" => DATA <= x"3036";
            when "01" & x"40a" => DATA <= x"3030";
            when "01" & x"40b" => DATA <= x"3730";
            when "01" & x"40c" => DATA <= x"3330";
            when "01" & x"40d" => DATA <= x"304b";
            when "01" & x"40e" => DATA <= x"070d";
            when "01" & x"40f" => DATA <= x"0a0d";
            when "01" & x"410" => DATA <= x"0a00";
            when "01" & x"411" => DATA <= x"1701";
            when "01" & x"412" => DATA <= x"0000";
            when "01" & x"413" => DATA <= x"0000";
            when "01" & x"414" => DATA <= x"0000";
            when "01" & x"415" => DATA <= x"0000";
            when "01" & x"416" => DATA <= x"0017";
            when "01" & x"417" => DATA <= x"0101";
            when "01" & x"418" => DATA <= x"0000";
            when "01" & x"419" => DATA <= x"0000";
            when "01" & x"41a" => DATA <= x"0000";
            when "01" & x"41b" => DATA <= x"0000";
            when "01" & x"41c" => DATA <= x"0a0d";
            when "01" & x"41d" => DATA <= x"4369";
            when "01" & x"41e" => DATA <= x"7363";
            when "01" & x"41f" => DATA <= x"4f53";
            when "01" & x"420" => DATA <= x"2076";
            when "01" & x"421" => DATA <= x"322e";
            when "01" & x"422" => DATA <= x"3031";
            when "01" & x"423" => DATA <= x"2028";
            when "01" & x"424" => DATA <= x"4a75";
            when "01" & x"425" => DATA <= x"6c79";
            when "01" & x"426" => DATA <= x"2033";
            when "01" & x"427" => DATA <= x"312c";
            when "01" & x"428" => DATA <= x"2032";
            when "01" & x"429" => DATA <= x"3031";
            when "01" & x"42a" => DATA <= x"3529";
            when "01" & x"42b" => DATA <= x"0a0d";
            when "01" & x"42c" => DATA <= x"0020";
            when "01" & x"42d" => DATA <= x"2020";
            when "01" & x"42e" => DATA <= x"5357";
            when "01" & x"42f" => DATA <= x"490a";
            when "01" & x"430" => DATA <= x"0d20";
            when "01" & x"431" => DATA <= x"2020";
            when "01" & x"432" => DATA <= x"5455";
            when "01" & x"433" => DATA <= x"4245";
            when "01" & x"434" => DATA <= x"0a0d";
            when "01" & x"435" => DATA <= x"0020";
            when "01" & x"436" => DATA <= x"2020";
            when "01" & x"437" => DATA <= x"4552";
            when "01" & x"438" => DATA <= x"524f";
            when "01" & x"439" => DATA <= x"5220";
            when "01" & x"43a" => DATA <= x"286e";
            when "01" & x"43b" => DATA <= x"756d";
            when "01" & x"43c" => DATA <= x"6265";
            when "01" & x"43d" => DATA <= x"7229";
            when "01" & x"43e" => DATA <= x"203c";
            when "01" & x"43f" => DATA <= x"6d65";
            when "01" & x"440" => DATA <= x"7373";
            when "01" & x"441" => DATA <= x"6167";
            when "01" & x"442" => DATA <= x"653e";
            when "01" & x"443" => DATA <= x"0a0d";
            when "01" & x"444" => DATA <= x"2020";
            when "01" & x"445" => DATA <= x"2046";
            when "01" & x"446" => DATA <= x"4c41";
            when "01" & x"447" => DATA <= x"5348";
            when "01" & x"448" => DATA <= x"203c";
            when "01" & x"449" => DATA <= x"6673";
            when "01" & x"44a" => DATA <= x"703e";
            when "01" & x"44b" => DATA <= x"0a0d";
            when "01" & x"44c" => DATA <= x"2020";
            when "01" & x"44d" => DATA <= x"2047";
            when "01" & x"44e" => DATA <= x"4f20";
            when "01" & x"44f" => DATA <= x"3c61";
            when "01" & x"450" => DATA <= x"6464";
            when "01" & x"451" => DATA <= x"723e";
            when "01" & x"452" => DATA <= x"0a0d";
            when "01" & x"453" => DATA <= x"2020";
            when "01" & x"454" => DATA <= x"204d";
            when "01" & x"455" => DATA <= x"4f4e";
            when "01" & x"456" => DATA <= x"0a0d";
            when "01" & x"457" => DATA <= x"2020";
            when "01" & x"458" => DATA <= x"2051";
            when "01" & x"459" => DATA <= x"5549";
            when "01" & x"45a" => DATA <= x"540a";
            when "01" & x"45b" => DATA <= x"0d20";
            when "01" & x"45c" => DATA <= x"2020";
            when "01" & x"45d" => DATA <= x"545a";
            when "01" & x"45e" => DATA <= x"4150";
            when "01" & x"45f" => DATA <= x"2028";
            when "01" & x"460" => DATA <= x"6164";
            when "01" & x"461" => DATA <= x"6472";
            when "01" & x"462" => DATA <= x"290a";
            when "01" & x"463" => DATA <= x"0d20";
            when "01" & x"464" => DATA <= x"2020";
            when "01" & x"465" => DATA <= x"5846";
            when "01" & x"466" => DATA <= x"4552";
            when "01" & x"467" => DATA <= x"203c";
            when "01" & x"468" => DATA <= x"696f";
            when "01" & x"469" => DATA <= x"2061";
            when "01" & x"46a" => DATA <= x"6464";
            when "01" & x"46b" => DATA <= x"722e";
            when "01" & x"46c" => DATA <= x"3e20";
            when "01" & x"46d" => DATA <= x"3c61";
            when "01" & x"46e" => DATA <= x"6464";
            when "01" & x"46f" => DATA <= x"723e";
            when "01" & x"470" => DATA <= x"203c";
            when "01" & x"471" => DATA <= x"6c65";
            when "01" & x"472" => DATA <= x"6e67";
            when "01" & x"473" => DATA <= x"7468";
            when "01" & x"474" => DATA <= x"3e20";
            when "01" & x"475" => DATA <= x"2852";
            when "01" & x"476" => DATA <= x"7c57";
            when "01" & x"477" => DATA <= x"2920";
            when "01" & x"478" => DATA <= x"2853";
            when "01" & x"479" => DATA <= x"7c4d";
            when "01" & x"47a" => DATA <= x"290a";
            when "01" & x"47b" => DATA <= x"0d00";
            when "01" & x"47c" => DATA <= x"5379";
            when "01" & x"47d" => DATA <= x"6e74";
            when "01" & x"47e" => DATA <= x"6178";
            when "01" & x"47f" => DATA <= x"3a20";
            when "01" & x"480" => DATA <= x"4552";
            when "01" & x"481" => DATA <= x"524f";
            when "01" & x"482" => DATA <= x"5220";
            when "01" & x"483" => DATA <= x"286e";
            when "01" & x"484" => DATA <= x"756d";
            when "01" & x"485" => DATA <= x"6265";
            when "01" & x"486" => DATA <= x"7229";
            when "01" & x"487" => DATA <= x"203c";
            when "01" & x"488" => DATA <= x"6d65";
            when "01" & x"489" => DATA <= x"7373";
            when "01" & x"48a" => DATA <= x"6167";
            when "01" & x"48b" => DATA <= x"653e";
            when "01" & x"48c" => DATA <= x"0a0d";
            when "01" & x"48d" => DATA <= x"0053";
            when "01" & x"48e" => DATA <= x"796e";
            when "01" & x"48f" => DATA <= x"7461";
            when "01" & x"490" => DATA <= x"783a";
            when "01" & x"491" => DATA <= x"2046";
            when "01" & x"492" => DATA <= x"4c41";
            when "01" & x"493" => DATA <= x"5348";
            when "01" & x"494" => DATA <= x"203c";
            when "01" & x"495" => DATA <= x"6673";
            when "01" & x"496" => DATA <= x"703e";
            when "01" & x"497" => DATA <= x"0a0d";
            when "01" & x"498" => DATA <= x"0053";
            when "01" & x"499" => DATA <= x"796e";
            when "01" & x"49a" => DATA <= x"7461";
            when "01" & x"49b" => DATA <= x"783a";
            when "01" & x"49c" => DATA <= x"2047";
            when "01" & x"49d" => DATA <= x"4f20";
            when "01" & x"49e" => DATA <= x"3c61";
            when "01" & x"49f" => DATA <= x"6464";
            when "01" & x"4a0" => DATA <= x"723e";
            when "01" & x"4a1" => DATA <= x"0a0d";
            when "01" & x"4a2" => DATA <= x"0053";
            when "01" & x"4a3" => DATA <= x"796e";
            when "01" & x"4a4" => DATA <= x"7461";
            when "01" & x"4a5" => DATA <= x"783a";
            when "01" & x"4a6" => DATA <= x"204d";
            when "01" & x"4a7" => DATA <= x"4f4e";
            when "01" & x"4a8" => DATA <= x"0a0d";
            when "01" & x"4a9" => DATA <= x"0053";
            when "01" & x"4aa" => DATA <= x"796e";
            when "01" & x"4ab" => DATA <= x"7461";
            when "01" & x"4ac" => DATA <= x"783a";
            when "01" & x"4ad" => DATA <= x"2054";
            when "01" & x"4ae" => DATA <= x"5a41";
            when "01" & x"4af" => DATA <= x"5020";
            when "01" & x"4b0" => DATA <= x"2861";
            when "01" & x"4b1" => DATA <= x"6464";
            when "01" & x"4b2" => DATA <= x"7229";
            when "01" & x"4b3" => DATA <= x"0a0d";
            when "01" & x"4b4" => DATA <= x"0053";
            when "01" & x"4b5" => DATA <= x"796e";
            when "01" & x"4b6" => DATA <= x"7461";
            when "01" & x"4b7" => DATA <= x"783a";
            when "01" & x"4b8" => DATA <= x"2058";
            when "01" & x"4b9" => DATA <= x"4645";
            when "01" & x"4ba" => DATA <= x"5220";
            when "01" & x"4bb" => DATA <= x"3c69";
            when "01" & x"4bc" => DATA <= x"6f20";
            when "01" & x"4bd" => DATA <= x"6164";
            when "01" & x"4be" => DATA <= x"6472";
            when "01" & x"4bf" => DATA <= x"2e3e";
            when "01" & x"4c0" => DATA <= x"203c";
            when "01" & x"4c1" => DATA <= x"6164";
            when "01" & x"4c2" => DATA <= x"6472";
            when "01" & x"4c3" => DATA <= x"3e20";
            when "01" & x"4c4" => DATA <= x"3c6c";
            when "01" & x"4c5" => DATA <= x"656e";
            when "01" & x"4c6" => DATA <= x"6774";
            when "01" & x"4c7" => DATA <= x"683e";
            when "01" & x"4c8" => DATA <= x"2028";
            when "01" & x"4c9" => DATA <= x"527c";
            when "01" & x"4ca" => DATA <= x"5729";
            when "01" & x"4cb" => DATA <= x"2028";
            when "01" & x"4cc" => DATA <= x"537c";
            when "01" & x"4cd" => DATA <= x"4d29";
            when "01" & x"4ce" => DATA <= x"0a0d";
            when "01" & x"4cf" => DATA <= x"0043";
            when "01" & x"4d0" => DATA <= x"6973";
            when "01" & x"4d1" => DATA <= x"634f";
            when "01" & x"4d2" => DATA <= x"5320";
            when "01" & x"4d3" => DATA <= x"4d6f";
            when "01" & x"4d4" => DATA <= x"6e69";
            when "01" & x"4d5" => DATA <= x"746f";
            when "01" & x"4d6" => DATA <= x"7200";
            when "01" & x"4d7" => DATA <= x"4220";
            when "01" & x"4d8" => DATA <= x"2042";
            when "01" & x"4d9" => DATA <= x"7974";
            when "01" & x"4da" => DATA <= x"6520";
            when "01" & x"4db" => DATA <= x"7365";
            when "01" & x"4dc" => DATA <= x"6172";
            when "01" & x"4dd" => DATA <= x"6368";
            when "01" & x"4de" => DATA <= x"203c";
            when "01" & x"4df" => DATA <= x"7374";
            when "01" & x"4e0" => DATA <= x"6172";
            when "01" & x"4e1" => DATA <= x"743e";
            when "01" & x"4e2" => DATA <= x"203c";
            when "01" & x"4e3" => DATA <= x"656e";
            when "01" & x"4e4" => DATA <= x"643e";
            when "01" & x"4e5" => DATA <= x"203c";
            when "01" & x"4e6" => DATA <= x"6279";
            when "01" & x"4e7" => DATA <= x"7465";
            when "01" & x"4e8" => DATA <= x"3e0a";
            when "01" & x"4e9" => DATA <= x"0d44";
            when "01" & x"4ea" => DATA <= x"2020";
            when "01" & x"4eb" => DATA <= x"4469";
            when "01" & x"4ec" => DATA <= x"7361";
            when "01" & x"4ed" => DATA <= x"7373";
            when "01" & x"4ee" => DATA <= x"656d";
            when "01" & x"4ef" => DATA <= x"626c";
            when "01" & x"4f0" => DATA <= x"6520";
            when "01" & x"4f1" => DATA <= x"3c61";
            when "01" & x"4f2" => DATA <= x"6464";
            when "01" & x"4f3" => DATA <= x"723e";
            when "01" & x"4f4" => DATA <= x"0a0d";
            when "01" & x"4f5" => DATA <= x"4520";
            when "01" & x"4f6" => DATA <= x"2045";
            when "01" & x"4f7" => DATA <= x"6469";
            when "01" & x"4f8" => DATA <= x"7420";
            when "01" & x"4f9" => DATA <= x"6d65";
            when "01" & x"4fa" => DATA <= x"6d6f";
            when "01" & x"4fb" => DATA <= x"7279";
            when "01" & x"4fc" => DATA <= x"203c";
            when "01" & x"4fd" => DATA <= x"6164";
            when "01" & x"4fe" => DATA <= x"6472";
            when "01" & x"4ff" => DATA <= x"3e0a";
            when "01" & x"500" => DATA <= x"0d46";
            when "01" & x"501" => DATA <= x"2020";
            when "01" & x"502" => DATA <= x"4669";
            when "01" & x"503" => DATA <= x"6c6c";
            when "01" & x"504" => DATA <= x"203c";
            when "01" & x"505" => DATA <= x"7374";
            when "01" & x"506" => DATA <= x"6172";
            when "01" & x"507" => DATA <= x"743e";
            when "01" & x"508" => DATA <= x"203c";
            when "01" & x"509" => DATA <= x"656e";
            when "01" & x"50a" => DATA <= x"643e";
            when "01" & x"50b" => DATA <= x"203c";
            when "01" & x"50c" => DATA <= x"6279";
            when "01" & x"50d" => DATA <= x"7465";
            when "01" & x"50e" => DATA <= x"3e0a";
            when "01" & x"50f" => DATA <= x"0d47";
            when "01" & x"510" => DATA <= x"2020";
            when "01" & x"511" => DATA <= x"476f";
            when "01" & x"512" => DATA <= x"203c";
            when "01" & x"513" => DATA <= x"6164";
            when "01" & x"514" => DATA <= x"6472";
            when "01" & x"515" => DATA <= x"3e0a";
            when "01" & x"516" => DATA <= x"0d48";
            when "01" & x"517" => DATA <= x"2020";
            when "01" & x"518" => DATA <= x"4865";
            when "01" & x"519" => DATA <= x"7820";
            when "01" & x"51a" => DATA <= x"6475";
            when "01" & x"51b" => DATA <= x"6d70";
            when "01" & x"51c" => DATA <= x"207b";
            when "01" & x"51d" => DATA <= x"6164";
            when "01" & x"51e" => DATA <= x"6472";
            when "01" & x"51f" => DATA <= x"7d0a";
            when "01" & x"520" => DATA <= x"0d4d";
            when "01" & x"521" => DATA <= x"2020";
            when "01" & x"522" => DATA <= x"4d6f";
            when "01" & x"523" => DATA <= x"7665";
            when "01" & x"524" => DATA <= x"206d";
            when "01" & x"525" => DATA <= x"656d";
            when "01" & x"526" => DATA <= x"6f72";
            when "01" & x"527" => DATA <= x"7920";
            when "01" & x"528" => DATA <= x"3c73";
            when "01" & x"529" => DATA <= x"6f75";
            when "01" & x"52a" => DATA <= x"7263";
            when "01" & x"52b" => DATA <= x"653e";
            when "01" & x"52c" => DATA <= x"203c";
            when "01" & x"52d" => DATA <= x"6465";
            when "01" & x"52e" => DATA <= x"7374";
            when "01" & x"52f" => DATA <= x"6e3e";
            when "01" & x"530" => DATA <= x"203c";
            when "01" & x"531" => DATA <= x"6c65";
            when "01" & x"532" => DATA <= x"6e67";
            when "01" & x"533" => DATA <= x"7468";
            when "01" & x"534" => DATA <= x"3e0a";
            when "01" & x"535" => DATA <= x"0d51";
            when "01" & x"536" => DATA <= x"2020";
            when "01" & x"537" => DATA <= x"5175";
            when "01" & x"538" => DATA <= x"6974";
            when "01" & x"539" => DATA <= x"0a0d";
            when "01" & x"53a" => DATA <= x"5220";
            when "01" & x"53b" => DATA <= x"2053";
            when "01" & x"53c" => DATA <= x"6574";
            when "01" & x"53d" => DATA <= x"2072";
            when "01" & x"53e" => DATA <= x"6567";
            when "01" & x"53f" => DATA <= x"6973";
            when "01" & x"540" => DATA <= x"7465";
            when "01" & x"541" => DATA <= x"7220";
            when "01" & x"542" => DATA <= x"636f";
            when "01" & x"543" => DATA <= x"6e74";
            when "01" & x"544" => DATA <= x"656e";
            when "01" & x"545" => DATA <= x"7473";
            when "01" & x"546" => DATA <= x"203c";
            when "01" & x"547" => DATA <= x"7265";
            when "01" & x"548" => DATA <= x"673e";
            when "01" & x"549" => DATA <= x"203c";
            when "01" & x"54a" => DATA <= x"7661";
            when "01" & x"54b" => DATA <= x"6c75";
            when "01" & x"54c" => DATA <= x"653e";
            when "01" & x"54d" => DATA <= x"0a0d";
            when "01" & x"54e" => DATA <= x"5320";
            when "01" & x"54f" => DATA <= x"2053";
            when "01" & x"550" => DATA <= x"7472";
            when "01" & x"551" => DATA <= x"696e";
            when "01" & x"552" => DATA <= x"6720";
            when "01" & x"553" => DATA <= x"7365";
            when "01" & x"554" => DATA <= x"6172";
            when "01" & x"555" => DATA <= x"6368";
            when "01" & x"556" => DATA <= x"203c";
            when "01" & x"557" => DATA <= x"7374";
            when "01" & x"558" => DATA <= x"6172";
            when "01" & x"559" => DATA <= x"743e";
            when "01" & x"55a" => DATA <= x"203c";
            when "01" & x"55b" => DATA <= x"656e";
            when "01" & x"55c" => DATA <= x"643e";
            when "01" & x"55d" => DATA <= x"203c";
            when "01" & x"55e" => DATA <= x"7374";
            when "01" & x"55f" => DATA <= x"7269";
            when "01" & x"560" => DATA <= x"6e67";
            when "01" & x"561" => DATA <= x"3e0a";
            when "01" & x"562" => DATA <= x"0d54";
            when "01" & x"563" => DATA <= x"2020";
            when "01" & x"564" => DATA <= x"5472";
            when "01" & x"565" => DATA <= x"6163";
            when "01" & x"566" => DATA <= x"650a";
            when "01" & x"567" => DATA <= x"0d56";
            when "01" & x"568" => DATA <= x"2020";
            when "01" & x"569" => DATA <= x"5669";
            when "01" & x"56a" => DATA <= x"6577";
            when "01" & x"56b" => DATA <= x"2072";
            when "01" & x"56c" => DATA <= x"6567";
            when "01" & x"56d" => DATA <= x"6973";
            when "01" & x"56e" => DATA <= x"7465";
            when "01" & x"56f" => DATA <= x"7220";
            when "01" & x"570" => DATA <= x"636f";
            when "01" & x"571" => DATA <= x"6e74";
            when "01" & x"572" => DATA <= x"656e";
            when "01" & x"573" => DATA <= x"7473";
            when "01" & x"574" => DATA <= x"0a0d";
            when "01" & x"575" => DATA <= x"2a20";
            when "01" & x"576" => DATA <= x"204f";
            when "01" & x"577" => DATA <= x"5320";
            when "01" & x"578" => DATA <= x"636f";
            when "01" & x"579" => DATA <= x"6d6d";
            when "01" & x"57a" => DATA <= x"616e";
            when "01" & x"57b" => DATA <= x"640a";
            when "01" & x"57c" => DATA <= x"0d3f";
            when "01" & x"57d" => DATA <= x"2020";
            when "01" & x"57e" => DATA <= x"4865";
            when "01" & x"57f" => DATA <= x"6c70";
            when "01" & x"580" => DATA <= x"0a0d";
            when "01" & x"581" => DATA <= x"0055";
            when "01" & x"582" => DATA <= x"6e6b";
            when "01" & x"583" => DATA <= x"6e6f";
            when "01" & x"584" => DATA <= x"776e";
            when "01" & x"585" => DATA <= x"2063";
            when "01" & x"586" => DATA <= x"6f6d";
            when "01" & x"587" => DATA <= x"6d61";
            when "01" & x"588" => DATA <= x"6e64";
            when "01" & x"589" => DATA <= x"2c20";
            when "01" & x"58a" => DATA <= x"7573";
            when "01" & x"58b" => DATA <= x"6520";
            when "01" & x"58c" => DATA <= x"3f20";
            when "01" & x"58d" => DATA <= x"666f";
            when "01" & x"58e" => DATA <= x"7220";
            when "01" & x"58f" => DATA <= x"6865";
            when "01" & x"590" => DATA <= x"6c70";
            when "01" & x"591" => DATA <= x"2e0a";
            when "01" & x"592" => DATA <= x"0d00";
            when "01" & x"593" => DATA <= x"542d";
            when "01" & x"594" => DATA <= x"532d";
            when "01" & x"595" => DATA <= x"2d49";
            when "01" & x"596" => DATA <= x"4e54";
            when "01" & x"597" => DATA <= x"2d2d";
            when "01" & x"598" => DATA <= x"2d58";
            when "01" & x"599" => DATA <= x"4e5a";
            when "01" & x"59a" => DATA <= x"5643";
            when "01" & x"59b" => DATA <= x"0046";
            when "01" & x"59c" => DATA <= x"696c";
            when "01" & x"59d" => DATA <= x"6520";
            when "01" & x"59e" => DATA <= x"6973";
            when "01" & x"59f" => DATA <= x"206e";
            when "01" & x"5a0" => DATA <= x"6f74";
            when "01" & x"5a1" => DATA <= x"2061";
            when "01" & x"5a2" => DATA <= x"2043";
            when "01" & x"5a3" => DATA <= x"6973";
            when "01" & x"5a4" => DATA <= x"634f";
            when "01" & x"5a5" => DATA <= x"5320";
            when "01" & x"5a6" => DATA <= x"6669";
            when "01" & x"5a7" => DATA <= x"6c65";
            when "01" & x"5a8" => DATA <= x"0a0d";
            when "01" & x"5a9" => DATA <= x"004e";
            when "01" & x"5aa" => DATA <= x"6f20";
            when "01" & x"5ab" => DATA <= x"726f";
            when "01" & x"5ac" => DATA <= x"6f6d";
            when "01" & x"5ad" => DATA <= x"0a0d";
            when "01" & x"5ae" => DATA <= x"0057";
            when "01" & x"5af" => DATA <= x"4152";
            when "01" & x"5b0" => DATA <= x"4e49";
            when "01" & x"5b1" => DATA <= x"4e47";
            when "01" & x"5b2" => DATA <= x"2120";
            when "01" & x"5b3" => DATA <= x"5448";
            when "01" & x"5b4" => DATA <= x"4953";
            when "01" & x"5b5" => DATA <= x"2057";
            when "01" & x"5b6" => DATA <= x"494c";
            when "01" & x"5b7" => DATA <= x"4c20";
            when "01" & x"5b8" => DATA <= x"464c";
            when "01" & x"5b9" => DATA <= x"4153";
            when "01" & x"5ba" => DATA <= x"4820";
            when "01" & x"5bb" => DATA <= x"5448";
            when "01" & x"5bc" => DATA <= x"4520";
            when "01" & x"5bd" => DATA <= x"4249";
            when "01" & x"5be" => DATA <= x"4f53";
            when "01" & x"5bf" => DATA <= x"0a0d";
            when "01" & x"5c0" => DATA <= x"5553";
            when "01" & x"5c1" => DATA <= x"4520";
            when "01" & x"5c2" => DATA <= x"4154";
            when "01" & x"5c3" => DATA <= x"2059";
            when "01" & x"5c4" => DATA <= x"4f55";
            when "01" & x"5c5" => DATA <= x"5220";
            when "01" & x"5c6" => DATA <= x"4f57";
            when "01" & x"5c7" => DATA <= x"4e20";
            when "01" & x"5c8" => DATA <= x"5249";
            when "01" & x"5c9" => DATA <= x"534b";
            when "01" & x"5ca" => DATA <= x"210a";
            when "01" & x"5cb" => DATA <= x"0d0a";
            when "01" & x"5cc" => DATA <= x"0d44";
            when "01" & x"5cd" => DATA <= x"6f20";
            when "01" & x"5ce" => DATA <= x"796f";
            when "01" & x"5cf" => DATA <= x"7520";
            when "01" & x"5d0" => DATA <= x"7761";
            when "01" & x"5d1" => DATA <= x"6e74";
            when "01" & x"5d2" => DATA <= x"2074";
            when "01" & x"5d3" => DATA <= x"6f20";
            when "01" & x"5d4" => DATA <= x"636f";
            when "01" & x"5d5" => DATA <= x"6e74";
            when "01" & x"5d6" => DATA <= x"696e";
            when "01" & x"5d7" => DATA <= x"7565";
            when "01" & x"5d8" => DATA <= x"3f20";
            when "01" & x"5d9" => DATA <= x"2859";
            when "01" & x"5da" => DATA <= x"2f4e";
            when "01" & x"5db" => DATA <= x"2920";
            when "01" & x"5dc" => DATA <= x"3a20";
            when "01" & x"5dd" => DATA <= x"0046";
            when "01" & x"5de" => DATA <= x"6c61";
            when "01" & x"5df" => DATA <= x"7368";
            when "01" & x"5e0" => DATA <= x"2052";
            when "01" & x"5e1" => DATA <= x"4f4d";
            when "01" & x"5e2" => DATA <= x"2049";
            when "01" & x"5e3" => DATA <= x"443d";
            when "01" & x"5e4" => DATA <= x"2400";
            when "01" & x"5e5" => DATA <= x"0a0d";
            when "01" & x"5e6" => DATA <= x"466c";
            when "01" & x"5e7" => DATA <= x"6173";
            when "01" & x"5e8" => DATA <= x"6869";
            when "01" & x"5e9" => DATA <= x"6e67";
            when "01" & x"5ea" => DATA <= x"2073";
            when "01" & x"5eb" => DATA <= x"6563";
            when "01" & x"5ec" => DATA <= x"746f";
            when "01" & x"5ed" => DATA <= x"7220";
            when "01" & x"5ee" => DATA <= x"0a0d";
            when "01" & x"5ef" => DATA <= x"0046";
            when "01" & x"5f0" => DATA <= x"6c61";
            when "01" & x"5f1" => DATA <= x"7368";
            when "01" & x"5f2" => DATA <= x"2063";
            when "01" & x"5f3" => DATA <= x"6f6d";
            when "01" & x"5f4" => DATA <= x"706c";
            when "01" & x"5f5" => DATA <= x"6574";
            when "01" & x"5f6" => DATA <= x"6564";
            when "01" & x"5f7" => DATA <= x"2073";
            when "01" & x"5f8" => DATA <= x"7563";
            when "01" & x"5f9" => DATA <= x"6365";
            when "01" & x"5fa" => DATA <= x"7373";
            when "01" & x"5fb" => DATA <= x"6675";
            when "01" & x"5fc" => DATA <= x"6c6c";
            when "01" & x"5fd" => DATA <= x"790a";
            when "01" & x"5fe" => DATA <= x"0d00";
            when "01" & x"5ff" => DATA <= x"466c";
            when "01" & x"600" => DATA <= x"6173";
            when "01" & x"601" => DATA <= x"6820";
            when "01" & x"602" => DATA <= x"6572";
            when "01" & x"603" => DATA <= x"726f";
            when "01" & x"604" => DATA <= x"7220";
            when "01" & x"605" => DATA <= x"6174";
            when "01" & x"606" => DATA <= x"2000";
            when "01" & x"607" => DATA <= x"4d6f";
            when "01" & x"608" => DATA <= x"6e54";
            when "01" & x"609" => DATA <= x"7565";
            when "01" & x"60a" => DATA <= x"5765";
            when "01" & x"60b" => DATA <= x"6454";
            when "01" & x"60c" => DATA <= x"6875";
            when "01" & x"60d" => DATA <= x"4672";
            when "01" & x"60e" => DATA <= x"6953";
            when "01" & x"60f" => DATA <= x"6174";
            when "01" & x"610" => DATA <= x"5375";
            when "01" & x"611" => DATA <= x"6e00";
            when "01" & x"612" => DATA <= x"4a61";
            when "01" & x"613" => DATA <= x"6e46";
            when "01" & x"614" => DATA <= x"6562";
            when "01" & x"615" => DATA <= x"4d61";
            when "01" & x"616" => DATA <= x"7241";
            when "01" & x"617" => DATA <= x"7072";
            when "01" & x"618" => DATA <= x"4d61";
            when "01" & x"619" => DATA <= x"794a";
            when "01" & x"61a" => DATA <= x"756e";
            when "01" & x"61b" => DATA <= x"4a75";
            when "01" & x"61c" => DATA <= x"6c41";
            when "01" & x"61d" => DATA <= x"7567";
            when "01" & x"61e" => DATA <= x"5365";
            when "01" & x"61f" => DATA <= x"704f";
            when "01" & x"620" => DATA <= x"6374";
            when "01" & x"621" => DATA <= x"4e6f";
            when "01" & x"622" => DATA <= x"7644";
            when "01" & x"623" => DATA <= x"6563";
            when "01" & x"624" => DATA <= x"000a";
            when "01" & x"625" => DATA <= x"0d42";
            when "01" & x"626" => DATA <= x"7573";
            when "01" & x"627" => DATA <= x"2065";
            when "01" & x"628" => DATA <= x"7272";
            when "01" & x"629" => DATA <= x"6f72";
            when "01" & x"62a" => DATA <= x"2061";
            when "01" & x"62b" => DATA <= x"7420";
            when "01" & x"62c" => DATA <= x"2400";
            when "01" & x"62d" => DATA <= x"0a0d";
            when "01" & x"62e" => DATA <= x"4164";
            when "01" & x"62f" => DATA <= x"6472";
            when "01" & x"630" => DATA <= x"6573";
            when "01" & x"631" => DATA <= x"7320";
            when "01" & x"632" => DATA <= x"6572";
            when "01" & x"633" => DATA <= x"726f";
            when "01" & x"634" => DATA <= x"7220";
            when "01" & x"635" => DATA <= x"6578";
            when "01" & x"636" => DATA <= x"6365";
            when "01" & x"637" => DATA <= x"7074";
            when "01" & x"638" => DATA <= x"696f";
            when "01" & x"639" => DATA <= x"6e20";
            when "01" & x"63a" => DATA <= x"6174";
            when "01" & x"63b" => DATA <= x"2024";
            when "01" & x"63c" => DATA <= x"0020";
            when "01" & x"63d" => DATA <= x"4163";
            when "01" & x"63e" => DATA <= x"6365";
            when "01" & x"63f" => DATA <= x"7373";
            when "01" & x"640" => DATA <= x"2074";
            when "01" & x"641" => DATA <= x"7970";
            when "01" & x"642" => DATA <= x"6526";
            when "01" & x"643" => DATA <= x"6675";
            when "01" & x"644" => DATA <= x"6e63";
            when "01" & x"645" => DATA <= x"7469";
            when "01" & x"646" => DATA <= x"6f6e";
            when "01" & x"647" => DATA <= x"3a00";
            when "01" & x"648" => DATA <= x"2041";
            when "01" & x"649" => DATA <= x"6363";
            when "01" & x"64a" => DATA <= x"6573";
            when "01" & x"64b" => DATA <= x"7320";
            when "01" & x"64c" => DATA <= x"6164";
            when "01" & x"64d" => DATA <= x"6472";
            when "01" & x"64e" => DATA <= x"6573";
            when "01" & x"64f" => DATA <= x"7320";
            when "01" & x"650" => DATA <= x"2020";
            when "01" & x"651" => DATA <= x"2020";
            when "01" & x"652" => DATA <= x"203a";
            when "01" & x"653" => DATA <= x"0020";
            when "01" & x"654" => DATA <= x"496e";
            when "01" & x"655" => DATA <= x"7374";
            when "01" & x"656" => DATA <= x"7275";
            when "01" & x"657" => DATA <= x"6374";
            when "01" & x"658" => DATA <= x"696f";
            when "01" & x"659" => DATA <= x"6e20";
            when "01" & x"65a" => DATA <= x"7265";
            when "01" & x"65b" => DATA <= x"6769";
            when "01" & x"65c" => DATA <= x"7374";
            when "01" & x"65d" => DATA <= x"6572";
            when "01" & x"65e" => DATA <= x"3a00";
            when "01" & x"65f" => DATA <= x"2053";
            when "01" & x"660" => DATA <= x"7461";
            when "01" & x"661" => DATA <= x"7475";
            when "01" & x"662" => DATA <= x"7320";
            when "01" & x"663" => DATA <= x"7265";
            when "01" & x"664" => DATA <= x"6769";
            when "01" & x"665" => DATA <= x"7374";
            when "01" & x"666" => DATA <= x"6572";
            when "01" & x"667" => DATA <= x"2020";
            when "01" & x"668" => DATA <= x"2020";
            when "01" & x"669" => DATA <= x"203a";
            when "01" & x"66a" => DATA <= x"5452";
            when "01" & x"66b" => DATA <= x"534d";
            when "01" & x"66c" => DATA <= x"2d49";
            when "01" & x"66d" => DATA <= x"4e54";
            when "01" & x"66e" => DATA <= x"2d2d";
            when "01" & x"66f" => DATA <= x"2d58";
            when "01" & x"670" => DATA <= x"4e5a";
            when "01" & x"671" => DATA <= x"5643";
            when "01" & x"672" => DATA <= x"0a0d";
            when "01" & x"673" => DATA <= x"2020";
            when "01" & x"674" => DATA <= x"2020";
            when "01" & x"675" => DATA <= x"2020";
            when "01" & x"676" => DATA <= x"2020";
            when "01" & x"677" => DATA <= x"2020";
            when "01" & x"678" => DATA <= x"2020";
            when "01" & x"679" => DATA <= x"2020";
            when "01" & x"67a" => DATA <= x"2020";
            when "01" & x"67b" => DATA <= x"2020";
            when "01" & x"67c" => DATA <= x"2020";
            when "01" & x"67d" => DATA <= x"2020";
            when "01" & x"67e" => DATA <= x"0000";
            when "01" & x"67f" => DATA <= x"0100";
            when "01" & x"680" => DATA <= x"8000";
            when "01" & x"681" => DATA <= x"0100";
            when "01" & x"682" => DATA <= x"496c";
            when "01" & x"683" => DATA <= x"6c65";
            when "01" & x"684" => DATA <= x"6761";
            when "01" & x"685" => DATA <= x"6c20";
            when "01" & x"686" => DATA <= x"696e";
            when "01" & x"687" => DATA <= x"7374";
            when "01" & x"688" => DATA <= x"7275";
            when "01" & x"689" => DATA <= x"6374";
            when "01" & x"68a" => DATA <= x"696f";
            when "01" & x"68b" => DATA <= x"6e00";
            when "01" & x"68c" => DATA <= x"8000";
            when "01" & x"68d" => DATA <= x"0104";
            when "01" & x"68e" => DATA <= x"556e";
            when "01" & x"68f" => DATA <= x"6b6e";
            when "01" & x"690" => DATA <= x"6f77";
            when "01" & x"691" => DATA <= x"6e20";
            when "01" & x"692" => DATA <= x"4952";
            when "01" & x"693" => DATA <= x"5120";
            when "01" & x"694" => DATA <= x"6174";
            when "01" & x"695" => DATA <= x"2026";
            when "01" & x"696" => DATA <= x"0000";
            when "01" & x"697" => DATA <= x"0169";
            when "01" & x"698" => DATA <= x"8000";
            when "01" & x"699" => DATA <= x"0169";
            when "01" & x"69a" => DATA <= x"496e";
            when "01" & x"69b" => DATA <= x"7465";
            when "01" & x"69c" => DATA <= x"6765";
            when "01" & x"69d" => DATA <= x"7220";
            when "01" & x"69e" => DATA <= x"6469";
            when "01" & x"69f" => DATA <= x"7669";
            when "01" & x"6a0" => DATA <= x"6465";
            when "01" & x"6a1" => DATA <= x"2062";
            when "01" & x"6a2" => DATA <= x"7920";
            when "01" & x"6a3" => DATA <= x"7a65";
            when "01" & x"6a4" => DATA <= x"726f";
            when "01" & x"6a5" => DATA <= x"0008";
            when "01" & x"6a6" => DATA <= x"8000";
            when "01" & x"6a7" => DATA <= x"0008";
            when "01" & x"6a8" => DATA <= x"5072";
            when "01" & x"6a9" => DATA <= x"6976";
            when "01" & x"6aa" => DATA <= x"696c";
            when "01" & x"6ab" => DATA <= x"6567";
            when "01" & x"6ac" => DATA <= x"6520";
            when "01" & x"6ad" => DATA <= x"7669";
            when "01" & x"6ae" => DATA <= x"6f6c";
            when "01" & x"6af" => DATA <= x"6174";
            when "01" & x"6b0" => DATA <= x"696f";
            when "01" & x"6b1" => DATA <= x"6e00";
            when "01" & x"6b2" => DATA <= x"0000";
            when "01" & x"6b3" => DATA <= x"0001";
            when "01" & x"6b4" => DATA <= x"4f75";
            when "01" & x"6b5" => DATA <= x"7420";
            when "01" & x"6b6" => DATA <= x"6f66";
            when "01" & x"6b7" => DATA <= x"2072";
            when "01" & x"6b8" => DATA <= x"616e";
            when "01" & x"6b9" => DATA <= x"6765";
            when "01" & x"6ba" => DATA <= x"0000";
            when "01" & x"6bb" => DATA <= x"0011";
            when "01" & x"6bc" => DATA <= x"0000";
            when "01" & x"6bd" => DATA <= x"0011";
            when "01" & x"6be" => DATA <= x"4573";
            when "01" & x"6bf" => DATA <= x"6361";
            when "01" & x"6c0" => DATA <= x"7065";
            when "01" & x"6c1" => DATA <= x"00ff";
            when "01" & x"6c2" => DATA <= x"0000";
            when "01" & x"6c3" => DATA <= x"00ff";
            when "01" & x"6c4" => DATA <= x"5468";
            when "01" & x"6c5" => DATA <= x"6973";
            when "01" & x"6c6" => DATA <= x"2069";
            when "01" & x"6c7" => DATA <= x"7320";
            when "01" & x"6c8" => DATA <= x"6e6f";
            when "01" & x"6c9" => DATA <= x"7420";
            when "01" & x"6ca" => DATA <= x"6120";
            when "01" & x"6cb" => DATA <= x"6c61";
            when "01" & x"6cc" => DATA <= x"6e67";
            when "01" & x"6cd" => DATA <= x"7561";
            when "01" & x"6ce" => DATA <= x"6765";
            when "01" & x"6cf" => DATA <= x"00ff";
            when "01" & x"6d0" => DATA <= x"0000";
            when "01" & x"6d1" => DATA <= x"00ff";
            when "01" & x"6d2" => DATA <= x"4920";
            when "01" & x"6d3" => DATA <= x"6361";
            when "01" & x"6d4" => DATA <= x"6e6e";
            when "01" & x"6d5" => DATA <= x"6f74";
            when "01" & x"6d6" => DATA <= x"2072";
            when "01" & x"6d7" => DATA <= x"756e";
            when "01" & x"6d8" => DATA <= x"2074";
            when "01" & x"6d9" => DATA <= x"6869";
            when "01" & x"6da" => DATA <= x"7320";
            when "01" & x"6db" => DATA <= x"636f";
            when "01" & x"6dc" => DATA <= x"6465";
            when "01" & x"6dd" => DATA <= x"00ff";
            when "01" & x"6de" => DATA <= x"0000";
            when "01" & x"6df" => DATA <= x"00ff";
            when "01" & x"6e0" => DATA <= x"556e";
            when "01" & x"6e1" => DATA <= x"6b6e";
            when "01" & x"6e2" => DATA <= x"6f77";
            when "01" & x"6e3" => DATA <= x"6e20";
            when "01" & x"6e4" => DATA <= x"6578";
            when "01" & x"6e5" => DATA <= x"6365";
            when "01" & x"6e6" => DATA <= x"7074";
            when "01" & x"6e7" => DATA <= x"696f";
            when "01" & x"6e8" => DATA <= x"6e00";
            when "01" & x"6e9" => DATA <= x"00ff";
            when "01" & x"6ea" => DATA <= x"0000";
            when "01" & x"6eb" => DATA <= x"00ff";
            when "01" & x"6ec" => DATA <= x"4e6f";
            when "01" & x"6ed" => DATA <= x"7420";
            when "01" & x"6ee" => DATA <= x"7375";
            when "01" & x"6ef" => DATA <= x"7070";
            when "01" & x"6f0" => DATA <= x"6f72";
            when "01" & x"6f1" => DATA <= x"7465";
            when "01" & x"6f2" => DATA <= x"6400";
            when "01" & x"6f3" => DATA <= x"016a";
            when "01" & x"6f4" => DATA <= x"0000";
            when "01" & x"6f5" => DATA <= x"016a";
            when "01" & x"6f6" => DATA <= x"4261";
            when "01" & x"6f7" => DATA <= x"6420";
            when "01" & x"6f8" => DATA <= x"6261";
            when "01" & x"6f9" => DATA <= x"7365";
            when "01" & x"6fa" => DATA <= x"0000";
            when "01" & x"6fb" => DATA <= x"016b";
            when "01" & x"6fc" => DATA <= x"0000";
            when "01" & x"6fd" => DATA <= x"016b";
            when "01" & x"6fe" => DATA <= x"4261";
            when "01" & x"6ff" => DATA <= x"6420";
            when "01" & x"700" => DATA <= x"6e75";
            when "01" & x"701" => DATA <= x"6d62";
            when "01" & x"702" => DATA <= x"6572";
            when "01" & x"703" => DATA <= x"006c";
            when "01" & x"704" => DATA <= x"0000";
            when "01" & x"705" => DATA <= x"016c";
            when "01" & x"706" => DATA <= x"4e75";
            when "01" & x"707" => DATA <= x"6d62";
            when "01" & x"708" => DATA <= x"6572";
            when "01" & x"709" => DATA <= x"2074";
            when "01" & x"70a" => DATA <= x"6f6f";
            when "01" & x"70b" => DATA <= x"2062";
            when "01" & x"70c" => DATA <= x"6967";
            when "01" & x"70d" => DATA <= x"00b0";
            when "01" & x"70e" => DATA <= x"0000";
            when "01" & x"70f" => DATA <= x"01b0";
            when "01" & x"710" => DATA <= x"4261";
            when "01" & x"711" => DATA <= x"6420";
            when "01" & x"712" => DATA <= x"656e";
            when "01" & x"713" => DATA <= x"7669";
            when "01" & x"714" => DATA <= x"726f";
            when "01" & x"715" => DATA <= x"6e6d";
            when "01" & x"716" => DATA <= x"656e";
            when "01" & x"717" => DATA <= x"7420";
            when "01" & x"718" => DATA <= x"6e75";
            when "01" & x"719" => DATA <= x"6d62";
            when "01" & x"71a" => DATA <= x"6572";
            when "01" & x"71b" => DATA <= x"00e6";
            when "01" & x"71c" => DATA <= x"0000";
            when "01" & x"71d" => DATA <= x"01e6";
            when "01" & x"71e" => DATA <= x"4e6f";
            when "01" & x"71f" => DATA <= x"2073";
            when "01" & x"720" => DATA <= x"7563";
            when "01" & x"721" => DATA <= x"6820";
            when "01" & x"722" => DATA <= x"5357";
            when "01" & x"723" => DATA <= x"4900";
            when "01" & x"724" => DATA <= x"0000";
            when "01" & x"725" => DATA <= x"01a0";
            when "01" & x"726" => DATA <= x"4261";
            when "01" & x"727" => DATA <= x"6420";
            when "01" & x"728" => DATA <= x"7665";
            when "01" & x"729" => DATA <= x"6374";
            when "01" & x"72a" => DATA <= x"6f72";
            when "01" & x"72b" => DATA <= x"206e";
            when "01" & x"72c" => DATA <= x"756d";
            when "01" & x"72d" => DATA <= x"6265";
            when "01" & x"72e" => DATA <= x"7200";
            when "01" & x"72f" => DATA <= x"01e2";
            when "01" & x"730" => DATA <= x"0000";
            when "01" & x"731" => DATA <= x"01e2";
            when "01" & x"732" => DATA <= x"5265";
            when "01" & x"733" => DATA <= x"7475";
            when "01" & x"734" => DATA <= x"726e";
            when "01" & x"735" => DATA <= x"2063";
            when "01" & x"736" => DATA <= x"6f64";
            when "01" & x"737" => DATA <= x"6520";
            when "01" & x"738" => DATA <= x"6c69";
            when "01" & x"739" => DATA <= x"6d69";
            when "01" & x"73a" => DATA <= x"7420";
            when "01" & x"73b" => DATA <= x"6578";
            when "01" & x"73c" => DATA <= x"6365";
            when "01" & x"73d" => DATA <= x"6564";
            when "01" & x"73e" => DATA <= x"6564";
            when "01" & x"73f" => DATA <= x"00e4";
            when "01" & x"740" => DATA <= x"0000";
            when "01" & x"741" => DATA <= x"01e4";
            when "01" & x"742" => DATA <= x"4275";
            when "01" & x"743" => DATA <= x"6666";
            when "01" & x"744" => DATA <= x"6572";
            when "01" & x"745" => DATA <= x"206f";
            when "01" & x"746" => DATA <= x"7665";
            when "01" & x"747" => DATA <= x"7266";
            when "01" & x"748" => DATA <= x"6c6f";
            when "01" & x"749" => DATA <= x"7700";
            when "01" & x"74a" => DATA <= x"0000";
            when "01" & x"74b" => DATA <= x"01e6";
            when "01" & x"74c" => DATA <= x"5357";
            when "01" & x"74d" => DATA <= x"4920";
            when "01" & x"74e" => DATA <= x"6e61";
            when "01" & x"74f" => DATA <= x"6d65";
            when "01" & x"750" => DATA <= x"206e";
            when "01" & x"751" => DATA <= x"6f74";
            when "01" & x"752" => DATA <= x"206b";
            when "01" & x"753" => DATA <= x"6e6f";
            when "01" & x"754" => DATA <= x"776e";
            when "01" & x"755" => DATA <= x"00c2";
            when "01" & x"756" => DATA <= x"0000";
            when "01" & x"757" => DATA <= x"02c2";
            when "01" & x"758" => DATA <= x"556e";
            when "01" & x"759" => DATA <= x"6b6e";
            when "01" & x"75a" => DATA <= x"6f77";
            when "01" & x"75b" => DATA <= x"6e20";
            when "01" & x"75c" => DATA <= x"2725";
            when "01" & x"75d" => DATA <= x"2720";
            when "01" & x"75e" => DATA <= x"6669";
            when "01" & x"75f" => DATA <= x"656c";
            when "01" & x"760" => DATA <= x"6400";
            when "01" & x"761" => DATA <= x"0306";
            when "01" & x"762" => DATA <= x"0000";
            when "01" & x"763" => DATA <= x"0306";
            when "01" & x"764" => DATA <= x"4261";
            when "01" & x"765" => DATA <= x"6420";
            when "01" & x"766" => DATA <= x"7374";
            when "01" & x"767" => DATA <= x"6174";
            when "01" & x"768" => DATA <= x"696f";
            when "01" & x"769" => DATA <= x"6e20";
            when "01" & x"76a" => DATA <= x"6e75";
            when "01" & x"76b" => DATA <= x"6d62";
            when "01" & x"76c" => DATA <= x"6572";
            when "01" & x"76d" => DATA <= x"0007";
            when "01" & x"76e" => DATA <= x"0000";
            when "01" & x"76f" => DATA <= x"0307";
            when "01" & x"770" => DATA <= x"4261";
            when "01" & x"771" => DATA <= x"6420";
            when "01" & x"772" => DATA <= x"6e65";
            when "01" & x"773" => DATA <= x"7477";
            when "01" & x"774" => DATA <= x"6f72";
            when "01" & x"775" => DATA <= x"6b20";
            when "01" & x"776" => DATA <= x"6e75";
            when "01" & x"777" => DATA <= x"6d62";
            when "01" & x"778" => DATA <= x"6572";
            when "01" & x"779" => DATA <= x"0001";
            when "01" & x"77a" => DATA <= x"0000";
            when "01" & x"77b" => DATA <= x"0401";
            when "01" & x"77c" => DATA <= x"4261";
            when "01" & x"77d" => DATA <= x"6420";
            when "01" & x"77e" => DATA <= x"4653";
            when "01" & x"77f" => DATA <= x"436f";
            when "01" & x"780" => DATA <= x"6e74";
            when "01" & x"781" => DATA <= x"726f";
            when "01" & x"782" => DATA <= x"6c20";
            when "01" & x"783" => DATA <= x"6361";
            when "01" & x"784" => DATA <= x"6c6c";
            when "01" & x"785" => DATA <= x"0007";
            when "01" & x"786" => DATA <= x"0000";
            when "01" & x"787" => DATA <= x"0807";
            when "01" & x"788" => DATA <= x"556e";
            when "01" & x"789" => DATA <= x"616c";
            when "01" & x"78a" => DATA <= x"6967";
            when "01" & x"78b" => DATA <= x"6e65";
            when "01" & x"78c" => DATA <= x"6420";
            when "01" & x"78d" => DATA <= x"6164";
            when "01" & x"78e" => DATA <= x"6472";
            when "01" & x"78f" => DATA <= x"6573";
            when "01" & x"790" => DATA <= x"7300";
            when "01" & x"791" => DATA <= x"0000";
            when "01" & x"792" => DATA <= x"0000";
            when "01" & x"793" => DATA <= x"0000";
            when "01" & x"794" => DATA <= x"0005";
            when "01" & x"795" => DATA <= x"0005";
            when "01" & x"796" => DATA <= x"0205";
            when "01" & x"797" => DATA <= x"080e";
            when "01" & x"798" => DATA <= x"0401";
            when "01" & x"799" => DATA <= x"0105";
            when "01" & x"79a" => DATA <= x"0001";
            when "01" & x"79b" => DATA <= x"2010";
            when "01" & x"79c" => DATA <= x"0d00";
            when "01" & x"79d" => DATA <= x"0480";
            when "01" & x"79e" => DATA <= x"0500";
            when "01" & x"79f" => DATA <= x"0500";
            when "01" & x"7a0" => DATA <= x"0500";
            when "01" & x"7a1" => DATA <= x"0000";
            when "01" & x"7a2" => DATA <= x"0509";
            when "01" & x"7a3" => DATA <= x"0500";
            when "01" & x"7a4" => DATA <= x"0818";
            when "01" & x"7a5" => DATA <= x"0001";
            when "01" & x"7a6" => DATA <= x"0d80";
            when "01" & x"7a7" => DATA <= x"0480";
            when "01" & x"7a8" => DATA <= x"0000";
            when "01" & x"7a9" => DATA <= x"0000";
            when "01" & x"7aa" => DATA <= x"003f";
            when "01" & x"7ab" => DATA <= x"09e6";
            when "01" & x"7ac" => DATA <= x"4f53";
            when "01" & x"7ad" => DATA <= x"5f57";
            when "01" & x"7ae" => DATA <= x"7269";
            when "01" & x"7af" => DATA <= x"7465";
            when "01" & x"7b0" => DATA <= x"4300";
            when "01" & x"7b1" => DATA <= x"0000";
            when "01" & x"7b2" => DATA <= x"0000";
            when "01" & x"7b3" => DATA <= x"0001";
            when "01" & x"7b4" => DATA <= x"003f";
            when "01" & x"7b5" => DATA <= x"09ec";
            when "01" & x"7b6" => DATA <= x"4f53";
            when "01" & x"7b7" => DATA <= x"5f57";
            when "01" & x"7b8" => DATA <= x"7269";
            when "01" & x"7b9" => DATA <= x"7465";
            when "01" & x"7ba" => DATA <= x"5300";
            when "01" & x"7bb" => DATA <= x"0000";
            when "01" & x"7bc" => DATA <= x"0000";
            when "01" & x"7bd" => DATA <= x"0002";
            when "01" & x"7be" => DATA <= x"003f";
            when "01" & x"7bf" => DATA <= x"09fe";
            when "01" & x"7c0" => DATA <= x"4f53";
            when "01" & x"7c1" => DATA <= x"5f57";
            when "01" & x"7c2" => DATA <= x"7269";
            when "01" & x"7c3" => DATA <= x"7465";
            when "01" & x"7c4" => DATA <= x"3000";
            when "01" & x"7c5" => DATA <= x"0000";
            when "01" & x"7c6" => DATA <= x"0000";
            when "01" & x"7c7" => DATA <= x"0003";
            when "01" & x"7c8" => DATA <= x"003f";
            when "01" & x"7c9" => DATA <= x"0a12";
            when "01" & x"7ca" => DATA <= x"4f53";
            when "01" & x"7cb" => DATA <= x"5f4e";
            when "01" & x"7cc" => DATA <= x"6577";
            when "01" & x"7cd" => DATA <= x"4c69";
            when "01" & x"7ce" => DATA <= x"6e65";
            when "01" & x"7cf" => DATA <= x"0000";
            when "01" & x"7d0" => DATA <= x"0000";
            when "01" & x"7d1" => DATA <= x"0004";
            when "01" & x"7d2" => DATA <= x"0000";
            when "01" & x"7d3" => DATA <= x"0410";
            when "01" & x"7d4" => DATA <= x"4f53";
            when "01" & x"7d5" => DATA <= x"5f52";
            when "01" & x"7d6" => DATA <= x"6561";
            when "01" & x"7d7" => DATA <= x"6443";
            when "01" & x"7d8" => DATA <= x"0000";
            when "01" & x"7d9" => DATA <= x"0000";
            when "01" & x"7da" => DATA <= x"0000";
            when "01" & x"7db" => DATA <= x"0005";
            when "01" & x"7dc" => DATA <= x"0000";
            when "01" & x"7dd" => DATA <= x"0414";
            when "01" & x"7de" => DATA <= x"4f53";
            when "01" & x"7df" => DATA <= x"5f43";
            when "01" & x"7e0" => DATA <= x"4c49";
            when "01" & x"7e1" => DATA <= x"0000";
            when "01" & x"7e2" => DATA <= x"0000";
            when "01" & x"7e3" => DATA <= x"0006";
            when "01" & x"7e4" => DATA <= x"0000";
            when "01" & x"7e5" => DATA <= x"0418";
            when "01" & x"7e6" => DATA <= x"4f53";
            when "01" & x"7e7" => DATA <= x"5f42";
            when "01" & x"7e8" => DATA <= x"7974";
            when "01" & x"7e9" => DATA <= x"6500";
            when "01" & x"7ea" => DATA <= x"0000";
            when "01" & x"7eb" => DATA <= x"0007";
            when "01" & x"7ec" => DATA <= x"0000";
            when "01" & x"7ed" => DATA <= x"041c";
            when "01" & x"7ee" => DATA <= x"4f53";
            when "01" & x"7ef" => DATA <= x"5f57";
            when "01" & x"7f0" => DATA <= x"6f72";
            when "01" & x"7f1" => DATA <= x"6400";
            when "01" & x"7f2" => DATA <= x"0000";
            when "01" & x"7f3" => DATA <= x"0008";
            when "01" & x"7f4" => DATA <= x"0000";
            when "01" & x"7f5" => DATA <= x"0420";
            when "01" & x"7f6" => DATA <= x"4f53";
            when "01" & x"7f7" => DATA <= x"5f46";
            when "01" & x"7f8" => DATA <= x"696c";
            when "01" & x"7f9" => DATA <= x"6500";
            when "01" & x"7fa" => DATA <= x"0000";
            when "01" & x"7fb" => DATA <= x"0009";
            when "01" & x"7fc" => DATA <= x"0000";
            when "01" & x"7fd" => DATA <= x"0424";
            when "01" & x"7fe" => DATA <= x"4f53";
            when "01" & x"7ff" => DATA <= x"5f41";
            when "01" & x"800" => DATA <= x"7267";
            when "01" & x"801" => DATA <= x"7300";
            when "01" & x"802" => DATA <= x"0000";
            when "01" & x"803" => DATA <= x"000a";
            when "01" & x"804" => DATA <= x"0000";
            when "01" & x"805" => DATA <= x"0428";
            when "01" & x"806" => DATA <= x"4f53";
            when "01" & x"807" => DATA <= x"5f42";
            when "01" & x"808" => DATA <= x"4765";
            when "01" & x"809" => DATA <= x"7400";
            when "01" & x"80a" => DATA <= x"0000";
            when "01" & x"80b" => DATA <= x"000b";
            when "01" & x"80c" => DATA <= x"0000";
            when "01" & x"80d" => DATA <= x"042c";
            when "01" & x"80e" => DATA <= x"4f53";
            when "01" & x"80f" => DATA <= x"5f42";
            when "01" & x"810" => DATA <= x"5075";
            when "01" & x"811" => DATA <= x"7400";
            when "01" & x"812" => DATA <= x"0000";
            when "01" & x"813" => DATA <= x"000c";
            when "01" & x"814" => DATA <= x"0000";
            when "01" & x"815" => DATA <= x"0430";
            when "01" & x"816" => DATA <= x"4f53";
            when "01" & x"817" => DATA <= x"5f47";
            when "01" & x"818" => DATA <= x"4250";
            when "01" & x"819" => DATA <= x"4200";
            when "01" & x"81a" => DATA <= x"0000";
            when "01" & x"81b" => DATA <= x"000d";
            when "01" & x"81c" => DATA <= x"0000";
            when "01" & x"81d" => DATA <= x"0434";
            when "01" & x"81e" => DATA <= x"4f53";
            when "01" & x"81f" => DATA <= x"5f46";
            when "01" & x"820" => DATA <= x"696e";
            when "01" & x"821" => DATA <= x"6400";
            when "01" & x"822" => DATA <= x"0000";
            when "01" & x"823" => DATA <= x"000e";
            when "01" & x"824" => DATA <= x"0000";
            when "01" & x"825" => DATA <= x"0438";
            when "01" & x"826" => DATA <= x"4f53";
            when "01" & x"827" => DATA <= x"5f52";
            when "01" & x"828" => DATA <= x"6561";
            when "01" & x"829" => DATA <= x"644c";
            when "01" & x"82a" => DATA <= x"696e";
            when "01" & x"82b" => DATA <= x"6500";
            when "01" & x"82c" => DATA <= x"0000";
            when "01" & x"82d" => DATA <= x"000f";
            when "01" & x"82e" => DATA <= x"003f";
            when "01" & x"82f" => DATA <= x"0df8";
            when "01" & x"830" => DATA <= x"4f53";
            when "01" & x"831" => DATA <= x"5f43";
            when "01" & x"832" => DATA <= x"6f6e";
            when "01" & x"833" => DATA <= x"7472";
            when "01" & x"834" => DATA <= x"6f6c";
            when "01" & x"835" => DATA <= x"0000";
            when "01" & x"836" => DATA <= x"0000";
            when "01" & x"837" => DATA <= x"0010";
            when "01" & x"838" => DATA <= x"003f";
            when "01" & x"839" => DATA <= x"0e30";
            when "01" & x"83a" => DATA <= x"4f53";
            when "01" & x"83b" => DATA <= x"5f47";
            when "01" & x"83c" => DATA <= x"6574";
            when "01" & x"83d" => DATA <= x"456e";
            when "01" & x"83e" => DATA <= x"7600";
            when "01" & x"83f" => DATA <= x"0000";
            when "01" & x"840" => DATA <= x"0000";
            when "01" & x"841" => DATA <= x"0011";
            when "01" & x"842" => DATA <= x"003f";
            when "01" & x"843" => DATA <= x"0e44";
            when "01" & x"844" => DATA <= x"4f53";
            when "01" & x"845" => DATA <= x"5f45";
            when "01" & x"846" => DATA <= x"7869";
            when "01" & x"847" => DATA <= x"7400";
            when "01" & x"848" => DATA <= x"0000";
            when "01" & x"849" => DATA <= x"0012";
            when "01" & x"84a" => DATA <= x"003f";
            when "01" & x"84b" => DATA <= x"0e4a";
            when "01" & x"84c" => DATA <= x"4f53";
            when "01" & x"84d" => DATA <= x"5f53";
            when "01" & x"84e" => DATA <= x"6574";
            when "01" & x"84f" => DATA <= x"456e";
            when "01" & x"850" => DATA <= x"7600";
            when "01" & x"851" => DATA <= x"0000";
            when "01" & x"852" => DATA <= x"0000";
            when "01" & x"853" => DATA <= x"0013";
            when "01" & x"854" => DATA <= x"003f";
            when "01" & x"855" => DATA <= x"0e9a";
            when "01" & x"856" => DATA <= x"4f53";
            when "01" & x"857" => DATA <= x"5f49";
            when "01" & x"858" => DATA <= x"6e74";
            when "01" & x"859" => DATA <= x"4f6e";
            when "01" & x"85a" => DATA <= x"0000";
            when "01" & x"85b" => DATA <= x"0000";
            when "01" & x"85c" => DATA <= x"0000";
            when "01" & x"85d" => DATA <= x"0014";
            when "01" & x"85e" => DATA <= x"003f";
            when "01" & x"85f" => DATA <= x"0ea0";
            when "01" & x"860" => DATA <= x"4f53";
            when "01" & x"861" => DATA <= x"5f49";
            when "01" & x"862" => DATA <= x"6e74";
            when "01" & x"863" => DATA <= x"4f66";
            when "01" & x"864" => DATA <= x"6600";
            when "01" & x"865" => DATA <= x"0000";
            when "01" & x"866" => DATA <= x"0000";
            when "01" & x"867" => DATA <= x"0015";
            when "01" & x"868" => DATA <= x"003f";
            when "01" & x"869" => DATA <= x"0ea6";
            when "01" & x"86a" => DATA <= x"4f53";
            when "01" & x"86b" => DATA <= x"5f43";
            when "01" & x"86c" => DATA <= x"616c";
            when "01" & x"86d" => DATA <= x"6c42";
            when "01" & x"86e" => DATA <= x"6163";
            when "01" & x"86f" => DATA <= x"6b00";
            when "01" & x"870" => DATA <= x"0000";
            when "01" & x"871" => DATA <= x"0016";
            when "01" & x"872" => DATA <= x"003f";
            when "01" & x"873" => DATA <= x"0ec6";
            when "01" & x"874" => DATA <= x"4f53";
            when "01" & x"875" => DATA <= x"5f45";
            when "01" & x"876" => DATA <= x"6e74";
            when "01" & x"877" => DATA <= x"6572";
            when "01" & x"878" => DATA <= x"4f53";
            when "01" & x"879" => DATA <= x"0000";
            when "01" & x"87a" => DATA <= x"0000";
            when "01" & x"87b" => DATA <= x"0018";
            when "01" & x"87c" => DATA <= x"003f";
            when "01" & x"87d" => DATA <= x"0ecc";
            when "01" & x"87e" => DATA <= x"4f53";
            when "01" & x"87f" => DATA <= x"5f42";
            when "01" & x"880" => DATA <= x"7265";
            when "01" & x"881" => DATA <= x"616b";
            when "01" & x"882" => DATA <= x"4374";
            when "01" & x"883" => DATA <= x"726c";
            when "01" & x"884" => DATA <= x"0000";
            when "01" & x"885" => DATA <= x"0000";
            when "01" & x"886" => DATA <= x"0000";
            when "01" & x"887" => DATA <= x"0019";
            when "01" & x"888" => DATA <= x"003f";
            when "01" & x"889" => DATA <= x"0eec";
            when "01" & x"88a" => DATA <= x"4f53";
            when "01" & x"88b" => DATA <= x"5f55";
            when "01" & x"88c" => DATA <= x"6e75";
            when "01" & x"88d" => DATA <= x"7365";
            when "01" & x"88e" => DATA <= x"6453";
            when "01" & x"88f" => DATA <= x"5749";
            when "01" & x"890" => DATA <= x"0000";
            when "01" & x"891" => DATA <= x"0000";
            when "01" & x"892" => DATA <= x"0000";
            when "01" & x"893" => DATA <= x"001c";
            when "01" & x"894" => DATA <= x"0000";
            when "01" & x"895" => DATA <= x"0468";
            when "01" & x"896" => DATA <= x"4f53";
            when "01" & x"897" => DATA <= x"5f4d";
            when "01" & x"898" => DATA <= x"6f75";
            when "01" & x"899" => DATA <= x"7365";
            when "01" & x"89a" => DATA <= x"0000";
            when "01" & x"89b" => DATA <= x"0000";
            when "01" & x"89c" => DATA <= x"0000";
            when "01" & x"89d" => DATA <= x"0021";
            when "01" & x"89e" => DATA <= x"003f";
            when "01" & x"89f" => DATA <= x"0fcc";
            when "01" & x"8a0" => DATA <= x"4f53";
            when "01" & x"8a1" => DATA <= x"5f52";
            when "01" & x"8a2" => DATA <= x"6561";
            when "01" & x"8a3" => DATA <= x"6455";
            when "01" & x"8a4" => DATA <= x"6e73";
            when "01" & x"8a5" => DATA <= x"6967";
            when "01" & x"8a6" => DATA <= x"6e65";
            when "01" & x"8a7" => DATA <= x"6400";
            when "01" & x"8a8" => DATA <= x"0000";
            when "01" & x"8a9" => DATA <= x"0028";
            when "01" & x"8aa" => DATA <= x"003f";
            when "01" & x"8ab" => DATA <= x"10c6";
            when "01" & x"8ac" => DATA <= x"4f53";
            when "01" & x"8ad" => DATA <= x"5f42";
            when "01" & x"8ae" => DATA <= x"696e";
            when "01" & x"8af" => DATA <= x"6172";
            when "01" & x"8b0" => DATA <= x"7954";
            when "01" & x"8b1" => DATA <= x"6f44";
            when "01" & x"8b2" => DATA <= x"6563";
            when "01" & x"8b3" => DATA <= x"696d";
            when "01" & x"8b4" => DATA <= x"616c";
            when "01" & x"8b5" => DATA <= x"0000";
            when "01" & x"8b6" => DATA <= x"0000";
            when "01" & x"8b7" => DATA <= x"0029";
            when "01" & x"8b8" => DATA <= x"0000";
            when "01" & x"8b9" => DATA <= x"043c";
            when "01" & x"8ba" => DATA <= x"4f53";
            when "01" & x"8bb" => DATA <= x"5f46";
            when "01" & x"8bc" => DATA <= x"5343";
            when "01" & x"8bd" => DATA <= x"6f6e";
            when "01" & x"8be" => DATA <= x"7472";
            when "01" & x"8bf" => DATA <= x"6f6c";
            when "01" & x"8c0" => DATA <= x"0000";
            when "01" & x"8c1" => DATA <= x"0000";
            when "01" & x"8c2" => DATA <= x"0000";
            when "01" & x"8c3" => DATA <= x"002b";
            when "01" & x"8c4" => DATA <= x"003f";
            when "01" & x"8c5" => DATA <= x"1120";
            when "01" & x"8c6" => DATA <= x"4f53";
            when "01" & x"8c7" => DATA <= x"5f47";
            when "01" & x"8c8" => DATA <= x"656e";
            when "01" & x"8c9" => DATA <= x"6572";
            when "01" & x"8ca" => DATA <= x"6174";
            when "01" & x"8cb" => DATA <= x"6545";
            when "01" & x"8cc" => DATA <= x"7272";
            when "01" & x"8cd" => DATA <= x"6f72";
            when "01" & x"8ce" => DATA <= x"0000";
            when "01" & x"8cf" => DATA <= x"0000";
            when "01" & x"8d0" => DATA <= x"0000";
            when "01" & x"8d1" => DATA <= x"002c";
            when "01" & x"8d2" => DATA <= x"003f";
            when "01" & x"8d3" => DATA <= x"1126";
            when "01" & x"8d4" => DATA <= x"4f53";
            when "01" & x"8d5" => DATA <= x"5f52";
            when "01" & x"8d6" => DATA <= x"6561";
            when "01" & x"8d7" => DATA <= x"6445";
            when "01" & x"8d8" => DATA <= x"7363";
            when "01" & x"8d9" => DATA <= x"6170";
            when "01" & x"8da" => DATA <= x"6553";
            when "01" & x"8db" => DATA <= x"7461";
            when "01" & x"8dc" => DATA <= x"7465";
            when "01" & x"8dd" => DATA <= x"0000";
            when "01" & x"8de" => DATA <= x"0000";
            when "01" & x"8df" => DATA <= x"002f";
            when "01" & x"8e0" => DATA <= x"003f";
            when "01" & x"8e1" => DATA <= x"113c";
            when "01" & x"8e2" => DATA <= x"4f53";
            when "01" & x"8e3" => DATA <= x"5f52";
            when "01" & x"8e4" => DATA <= x"6561";
            when "01" & x"8e5" => DATA <= x"6450";
            when "01" & x"8e6" => DATA <= x"616c";
            when "01" & x"8e7" => DATA <= x"6574";
            when "01" & x"8e8" => DATA <= x"7465";
            when "01" & x"8e9" => DATA <= x"0000";
            when "01" & x"8ea" => DATA <= x"0000";
            when "01" & x"8eb" => DATA <= x"0032";
            when "01" & x"8ec" => DATA <= x"003f";
            when "01" & x"8ed" => DATA <= x"1152";
            when "01" & x"8ee" => DATA <= x"4f53";
            when "01" & x"8ef" => DATA <= x"5f52";
            when "01" & x"8f0" => DATA <= x"6561";
            when "01" & x"8f1" => DATA <= x"6450";
            when "01" & x"8f2" => DATA <= x"6f69";
            when "01" & x"8f3" => DATA <= x"6e74";
            when "01" & x"8f4" => DATA <= x"0000";
            when "01" & x"8f5" => DATA <= x"0000";
            when "01" & x"8f6" => DATA <= x"0000";
            when "01" & x"8f7" => DATA <= x"0034";
            when "01" & x"8f8" => DATA <= x"003f";
            when "01" & x"8f9" => DATA <= x"11a8";
            when "01" & x"8fa" => DATA <= x"4f53";
            when "01" & x"8fb" => DATA <= x"5f43";
            when "01" & x"8fc" => DATA <= x"616c";
            when "01" & x"8fd" => DATA <= x"6c41";
            when "01" & x"8fe" => DATA <= x"5665";
            when "01" & x"8ff" => DATA <= x"6374";
            when "01" & x"900" => DATA <= x"6f72";
            when "01" & x"901" => DATA <= x"0000";
            when "01" & x"902" => DATA <= x"0000";
            when "01" & x"903" => DATA <= x"0036";
            when "01" & x"904" => DATA <= x"003f";
            when "01" & x"905" => DATA <= x"11d4";
            when "01" & x"906" => DATA <= x"4f53";
            when "01" & x"907" => DATA <= x"5f52";
            when "01" & x"908" => DATA <= x"656d";
            when "01" & x"909" => DATA <= x"6f76";
            when "01" & x"90a" => DATA <= x"6543";
            when "01" & x"90b" => DATA <= x"7572";
            when "01" & x"90c" => DATA <= x"736f";
            when "01" & x"90d" => DATA <= x"7273";
            when "01" & x"90e" => DATA <= x"0000";
            when "01" & x"90f" => DATA <= x"0000";
            when "01" & x"910" => DATA <= x"0000";
            when "01" & x"911" => DATA <= x"0037";
            when "01" & x"912" => DATA <= x"003f";
            when "01" & x"913" => DATA <= x"11ee";
            when "01" & x"914" => DATA <= x"4f53";
            when "01" & x"915" => DATA <= x"5f52";
            when "01" & x"916" => DATA <= x"6573";
            when "01" & x"917" => DATA <= x"746f";
            when "01" & x"918" => DATA <= x"7265";
            when "01" & x"919" => DATA <= x"4375";
            when "01" & x"91a" => DATA <= x"7273";
            when "01" & x"91b" => DATA <= x"6f72";
            when "01" & x"91c" => DATA <= x"7300";
            when "01" & x"91d" => DATA <= x"0000";
            when "01" & x"91e" => DATA <= x"0000";
            when "01" & x"91f" => DATA <= x"0038";
            when "01" & x"920" => DATA <= x"003f";
            when "01" & x"921" => DATA <= x"1208";
            when "01" & x"922" => DATA <= x"4f53";
            when "01" & x"923" => DATA <= x"5f53";
            when "01" & x"924" => DATA <= x"5749";
            when "01" & x"925" => DATA <= x"4e75";
            when "01" & x"926" => DATA <= x"6d62";
            when "01" & x"927" => DATA <= x"6572";
            when "01" & x"928" => DATA <= x"546f";
            when "01" & x"929" => DATA <= x"5374";
            when "01" & x"92a" => DATA <= x"7269";
            when "01" & x"92b" => DATA <= x"6e67";
            when "01" & x"92c" => DATA <= x"0000";
            when "01" & x"92d" => DATA <= x"0000";
            when "01" & x"92e" => DATA <= x"0000";
            when "01" & x"92f" => DATA <= x"0039";
            when "01" & x"930" => DATA <= x"003f";
            when "01" & x"931" => DATA <= x"1288";
            when "01" & x"932" => DATA <= x"4f53";
            when "01" & x"933" => DATA <= x"5f53";
            when "01" & x"934" => DATA <= x"5749";
            when "01" & x"935" => DATA <= x"4e75";
            when "01" & x"936" => DATA <= x"6d62";
            when "01" & x"937" => DATA <= x"6572";
            when "01" & x"938" => DATA <= x"4672";
            when "01" & x"939" => DATA <= x"6f6d";
            when "01" & x"93a" => DATA <= x"5374";
            when "01" & x"93b" => DATA <= x"7269";
            when "01" & x"93c" => DATA <= x"6e67";
            when "01" & x"93d" => DATA <= x"0000";
            when "01" & x"93e" => DATA <= x"0000";
            when "01" & x"93f" => DATA <= x"003a";
            when "01" & x"940" => DATA <= x"003f";
            when "01" & x"941" => DATA <= x"12cc";
            when "01" & x"942" => DATA <= x"4f53";
            when "01" & x"943" => DATA <= x"5f56";
            when "01" & x"944" => DATA <= x"616c";
            when "01" & x"945" => DATA <= x"6964";
            when "01" & x"946" => DATA <= x"6174";
            when "01" & x"947" => DATA <= x"6541";
            when "01" & x"948" => DATA <= x"6464";
            when "01" & x"949" => DATA <= x"7265";
            when "01" & x"94a" => DATA <= x"7373";
            when "01" & x"94b" => DATA <= x"0000";
            when "01" & x"94c" => DATA <= x"0000";
            when "01" & x"94d" => DATA <= x"003f";
            when "01" & x"94e" => DATA <= x"003f";
            when "01" & x"94f" => DATA <= x"12e6";
            when "01" & x"950" => DATA <= x"4f53";
            when "01" & x"951" => DATA <= x"5f43";
            when "01" & x"952" => DATA <= x"6865";
            when "01" & x"953" => DATA <= x"636b";
            when "01" & x"954" => DATA <= x"4d6f";
            when "01" & x"955" => DATA <= x"6465";
            when "01" & x"956" => DATA <= x"5661";
            when "01" & x"957" => DATA <= x"6c69";
            when "01" & x"958" => DATA <= x"6400";
            when "01" & x"959" => DATA <= x"0000";
            when "01" & x"95a" => DATA <= x"0000";
            when "01" & x"95b" => DATA <= x"0040";
            when "01" & x"95c" => DATA <= x"003f";
            when "01" & x"95d" => DATA <= x"1300";
            when "01" & x"95e" => DATA <= x"4f53";
            when "01" & x"95f" => DATA <= x"5f43";
            when "01" & x"960" => DATA <= x"6861";
            when "01" & x"961" => DATA <= x"6e67";
            when "01" & x"962" => DATA <= x"6545";
            when "01" & x"963" => DATA <= x"6e76";
            when "01" & x"964" => DATA <= x"6972";
            when "01" & x"965" => DATA <= x"6f6e";
            when "01" & x"966" => DATA <= x"6d65";
            when "01" & x"967" => DATA <= x"6e74";
            when "01" & x"968" => DATA <= x"0000";
            when "01" & x"969" => DATA <= x"0000";
            when "01" & x"96a" => DATA <= x"0000";
            when "01" & x"96b" => DATA <= x"0042";
            when "01" & x"96c" => DATA <= x"003f";
            when "01" & x"96d" => DATA <= x"1306";
            when "01" & x"96e" => DATA <= x"4f53";
            when "01" & x"96f" => DATA <= x"5f52";
            when "01" & x"970" => DATA <= x"6561";
            when "01" & x"971" => DATA <= x"644d";
            when "01" & x"972" => DATA <= x"6f6e";
            when "01" & x"973" => DATA <= x"6f74";
            when "01" & x"974" => DATA <= x"6f6e";
            when "01" & x"975" => DATA <= x"6963";
            when "01" & x"976" => DATA <= x"5469";
            when "01" & x"977" => DATA <= x"6d65";
            when "01" & x"978" => DATA <= x"0000";
            when "01" & x"979" => DATA <= x"0000";
            when "01" & x"97a" => DATA <= x"0000";
            when "01" & x"97b" => DATA <= x"0045";
            when "01" & x"97c" => DATA <= x"003f";
            when "01" & x"97d" => DATA <= x"1320";
            when "01" & x"97e" => DATA <= x"4f53";
            when "01" & x"97f" => DATA <= x"5f50";
            when "01" & x"980" => DATA <= x"6c6f";
            when "01" & x"981" => DATA <= x"7400";
            when "01" & x"982" => DATA <= x"0000";
            when "01" & x"983" => DATA <= x"0046";
            when "01" & x"984" => DATA <= x"003f";
            when "01" & x"985" => DATA <= x"136e";
            when "01" & x"986" => DATA <= x"4f53";
            when "01" & x"987" => DATA <= x"5f57";
            when "01" & x"988" => DATA <= x"7269";
            when "01" & x"989" => DATA <= x"7465";
            when "01" & x"98a" => DATA <= x"4e00";
            when "01" & x"98b" => DATA <= x"0000";
            when "01" & x"98c" => DATA <= x"0000";
            when "01" & x"98d" => DATA <= x"0048";
            when "01" & x"98e" => DATA <= x"003f";
            when "01" & x"98f" => DATA <= x"1394";
            when "01" & x"990" => DATA <= x"4f53";
            when "01" & x"991" => DATA <= x"5f57";
            when "01" & x"992" => DATA <= x"7269";
            when "01" & x"993" => DATA <= x"7465";
            when "01" & x"994" => DATA <= x"456e";
            when "01" & x"995" => DATA <= x"7600";
            when "01" & x"996" => DATA <= x"0000";
            when "01" & x"997" => DATA <= x"0050";
            when "01" & x"998" => DATA <= x"003f";
            when "01" & x"999" => DATA <= x"13ca";
            when "01" & x"99a" => DATA <= x"4f53";
            when "01" & x"99b" => DATA <= x"5f45";
            when "01" & x"99c" => DATA <= x"7869";
            when "01" & x"99d" => DATA <= x"7441";
            when "01" & x"99e" => DATA <= x"6e64";
            when "01" & x"99f" => DATA <= x"4469";
            when "01" & x"9a0" => DATA <= x"6500";
            when "01" & x"9a1" => DATA <= x"0000";
            when "01" & x"9a2" => DATA <= x"0000";
            when "01" & x"9a3" => DATA <= x"0055";
            when "01" & x"9a4" => DATA <= x"003f";
            when "01" & x"9a5" => DATA <= x"13e2";
            when "01" & x"9a6" => DATA <= x"4f53";
            when "01" & x"9a7" => DATA <= x"5f52";
            when "01" & x"9a8" => DATA <= x"6561";
            when "01" & x"9a9" => DATA <= x"6444";
            when "01" & x"9aa" => DATA <= x"6566";
            when "01" & x"9ab" => DATA <= x"6175";
            when "01" & x"9ac" => DATA <= x"6c74";
            when "01" & x"9ad" => DATA <= x"4861";
            when "01" & x"9ae" => DATA <= x"6e64";
            when "01" & x"9af" => DATA <= x"6c65";
            when "01" & x"9b0" => DATA <= x"7200";
            when "01" & x"9b1" => DATA <= x"0000";
            when "01" & x"9b2" => DATA <= x"0000";
            when "01" & x"9b3" => DATA <= x"0056";
            when "01" & x"9b4" => DATA <= x"003f";
            when "01" & x"9b5" => DATA <= x"142a";
            when "01" & x"9b6" => DATA <= x"4f53";
            when "01" & x"9b7" => DATA <= x"5f53";
            when "01" & x"9b8" => DATA <= x"6574";
            when "01" & x"9b9" => DATA <= x"4543";
            when "01" & x"9ba" => DATA <= x"464f";
            when "01" & x"9bb" => DATA <= x"7269";
            when "01" & x"9bc" => DATA <= x"6769";
            when "01" & x"9bd" => DATA <= x"6e00";
            when "01" & x"9be" => DATA <= x"0000";
            when "01" & x"9bf" => DATA <= x"005d";
            when "01" & x"9c0" => DATA <= x"003f";
            when "01" & x"9c1" => DATA <= x"14da";
            when "01" & x"9c2" => DATA <= x"4f53";
            when "01" & x"9c3" => DATA <= x"5f50";
            when "01" & x"9c4" => DATA <= x"7269";
            when "01" & x"9c5" => DATA <= x"6e74";
            when "01" & x"9c6" => DATA <= x"4368";
            when "01" & x"9c7" => DATA <= x"6172";
            when "01" & x"9c8" => DATA <= x"0000";
            when "01" & x"9c9" => DATA <= x"0000";
            when "01" & x"9ca" => DATA <= x"0000";
            when "01" & x"9cb" => DATA <= x"005b";
            when "01" & x"9cc" => DATA <= x"003f";
            when "01" & x"9cd" => DATA <= x"14a8";
            when "01" & x"9ce" => DATA <= x"4f53";
            when "01" & x"9cf" => DATA <= x"5f43";
            when "01" & x"9d0" => DATA <= x"5243";
            when "01" & x"9d1" => DATA <= x"0000";
            when "01" & x"9d2" => DATA <= x"0000";
            when "01" & x"9d3" => DATA <= x"0059";
            when "01" & x"9d4" => DATA <= x"003f";
            when "01" & x"9d5" => DATA <= x"149a";
            when "01" & x"9d6" => DATA <= x"4f53";
            when "01" & x"9d7" => DATA <= x"5f43";
            when "01" & x"9d8" => DATA <= x"6f6e";
            when "01" & x"9d9" => DATA <= x"6669";
            when "01" & x"9da" => DATA <= x"726d";
            when "01" & x"9db" => DATA <= x"0000";
            when "01" & x"9dc" => DATA <= x"0000";
            when "01" & x"9dd" => DATA <= x"007c";
            when "01" & x"9de" => DATA <= x"003f";
            when "01" & x"9df" => DATA <= x"14e6";
            when "01" & x"9e0" => DATA <= x"4f53";
            when "01" & x"9e1" => DATA <= x"5f4c";
            when "01" & x"9e2" => DATA <= x"6561";
            when "01" & x"9e3" => DATA <= x"7665";
            when "01" & x"9e4" => DATA <= x"4f53";
            when "01" & x"9e5" => DATA <= x"0000";
            when "01" & x"9e6" => DATA <= x"0000";
            when "01" & x"9e7" => DATA <= x"007d";
            when "01" & x"9e8" => DATA <= x"003f";
            when "01" & x"9e9" => DATA <= x"14ec";
            when "01" & x"9ea" => DATA <= x"4f53";
            when "01" & x"9eb" => DATA <= x"5f52";
            when "01" & x"9ec" => DATA <= x"6561";
            when "01" & x"9ed" => DATA <= x"644c";
            when "01" & x"9ee" => DATA <= x"696e";
            when "01" & x"9ef" => DATA <= x"6533";
            when "01" & x"9f0" => DATA <= x"3200";
            when "01" & x"9f1" => DATA <= x"0000";
            when "01" & x"9f2" => DATA <= x"0000";
            when "01" & x"9f3" => DATA <= x"00d0";
            when "01" & x"9f4" => DATA <= x"003f";
            when "01" & x"9f5" => DATA <= x"1674";
            when "01" & x"9f6" => DATA <= x"4f53";
            when "01" & x"9f7" => DATA <= x"5f43";
            when "01" & x"9f8" => DATA <= x"6f6e";
            when "01" & x"9f9" => DATA <= x"7665";
            when "01" & x"9fa" => DATA <= x"7274";
            when "01" & x"9fb" => DATA <= x"4865";
            when "01" & x"9fc" => DATA <= x"7831";
            when "01" & x"9fd" => DATA <= x"0000";
            when "01" & x"9fe" => DATA <= x"0000";
            when "01" & x"9ff" => DATA <= x"00d1";
            when "01" & x"a00" => DATA <= x"003f";
            when "01" & x"a01" => DATA <= x"1690";
            when "01" & x"a02" => DATA <= x"4f53";
            when "01" & x"a03" => DATA <= x"5f43";
            when "01" & x"a04" => DATA <= x"6f6e";
            when "01" & x"a05" => DATA <= x"7665";
            when "01" & x"a06" => DATA <= x"7274";
            when "01" & x"a07" => DATA <= x"4865";
            when "01" & x"a08" => DATA <= x"7832";
            when "01" & x"a09" => DATA <= x"0000";
            when "01" & x"a0a" => DATA <= x"0000";
            when "01" & x"a0b" => DATA <= x"00d2";
            when "01" & x"a0c" => DATA <= x"003f";
            when "01" & x"a0d" => DATA <= x"16ac";
            when "01" & x"a0e" => DATA <= x"4f53";
            when "01" & x"a0f" => DATA <= x"5f43";
            when "01" & x"a10" => DATA <= x"6f6e";
            when "01" & x"a11" => DATA <= x"7665";
            when "01" & x"a12" => DATA <= x"7274";
            when "01" & x"a13" => DATA <= x"4865";
            when "01" & x"a14" => DATA <= x"7834";
            when "01" & x"a15" => DATA <= x"0000";
            when "01" & x"a16" => DATA <= x"0000";
            when "01" & x"a17" => DATA <= x"00d3";
            when "01" & x"a18" => DATA <= x"003f";
            when "01" & x"a19" => DATA <= x"16ca";
            when "01" & x"a1a" => DATA <= x"4f53";
            when "01" & x"a1b" => DATA <= x"5f43";
            when "01" & x"a1c" => DATA <= x"6f6e";
            when "01" & x"a1d" => DATA <= x"7665";
            when "01" & x"a1e" => DATA <= x"7274";
            when "01" & x"a1f" => DATA <= x"4865";
            when "01" & x"a20" => DATA <= x"7836";
            when "01" & x"a21" => DATA <= x"0000";
            when "01" & x"a22" => DATA <= x"0000";
            when "01" & x"a23" => DATA <= x"00d4";
            when "01" & x"a24" => DATA <= x"003f";
            when "01" & x"a25" => DATA <= x"16e6";
            when "01" & x"a26" => DATA <= x"4f53";
            when "01" & x"a27" => DATA <= x"5f43";
            when "01" & x"a28" => DATA <= x"6f6e";
            when "01" & x"a29" => DATA <= x"7665";
            when "01" & x"a2a" => DATA <= x"7274";
            when "01" & x"a2b" => DATA <= x"4865";
            when "01" & x"a2c" => DATA <= x"7838";
            when "01" & x"a2d" => DATA <= x"0000";
            when "01" & x"a2e" => DATA <= x"0000";
            when "01" & x"a2f" => DATA <= x"00d5";
            when "01" & x"a30" => DATA <= x"003f";
            when "01" & x"a31" => DATA <= x"1740";
            when "01" & x"a32" => DATA <= x"4f53";
            when "01" & x"a33" => DATA <= x"5f43";
            when "01" & x"a34" => DATA <= x"6f6e";
            when "01" & x"a35" => DATA <= x"7665";
            when "01" & x"a36" => DATA <= x"7274";
            when "01" & x"a37" => DATA <= x"4361";
            when "01" & x"a38" => DATA <= x"7264";
            when "01" & x"a39" => DATA <= x"696e";
            when "01" & x"a3a" => DATA <= x"616c";
            when "01" & x"a3b" => DATA <= x"3100";
            when "01" & x"a3c" => DATA <= x"0000";
            when "01" & x"a3d" => DATA <= x"00d6";
            when "01" & x"a3e" => DATA <= x"003f";
            when "01" & x"a3f" => DATA <= x"175a";
            when "01" & x"a40" => DATA <= x"4f53";
            when "01" & x"a41" => DATA <= x"5f43";
            when "01" & x"a42" => DATA <= x"6f6e";
            when "01" & x"a43" => DATA <= x"7665";
            when "01" & x"a44" => DATA <= x"7274";
            when "01" & x"a45" => DATA <= x"4361";
            when "01" & x"a46" => DATA <= x"7264";
            when "01" & x"a47" => DATA <= x"696e";
            when "01" & x"a48" => DATA <= x"616c";
            when "01" & x"a49" => DATA <= x"3200";
            when "01" & x"a4a" => DATA <= x"0000";
            when "01" & x"a4b" => DATA <= x"00d7";
            when "01" & x"a4c" => DATA <= x"003f";
            when "01" & x"a4d" => DATA <= x"1774";
            when "01" & x"a4e" => DATA <= x"4f53";
            when "01" & x"a4f" => DATA <= x"5f43";
            when "01" & x"a50" => DATA <= x"6f6e";
            when "01" & x"a51" => DATA <= x"7665";
            when "01" & x"a52" => DATA <= x"7274";
            when "01" & x"a53" => DATA <= x"4361";
            when "01" & x"a54" => DATA <= x"7264";
            when "01" & x"a55" => DATA <= x"696e";
            when "01" & x"a56" => DATA <= x"616c";
            when "01" & x"a57" => DATA <= x"3300";
            when "01" & x"a58" => DATA <= x"0000";
            when "01" & x"a59" => DATA <= x"00d8";
            when "01" & x"a5a" => DATA <= x"003f";
            when "01" & x"a5b" => DATA <= x"178e";
            when "01" & x"a5c" => DATA <= x"4f53";
            when "01" & x"a5d" => DATA <= x"5f43";
            when "01" & x"a5e" => DATA <= x"6f6e";
            when "01" & x"a5f" => DATA <= x"7665";
            when "01" & x"a60" => DATA <= x"7274";
            when "01" & x"a61" => DATA <= x"4361";
            when "01" & x"a62" => DATA <= x"7264";
            when "01" & x"a63" => DATA <= x"696e";
            when "01" & x"a64" => DATA <= x"616c";
            when "01" & x"a65" => DATA <= x"3400";
            when "01" & x"a66" => DATA <= x"0000";
            when "01" & x"a67" => DATA <= x"00d9";
            when "01" & x"a68" => DATA <= x"003f";
            when "01" & x"a69" => DATA <= x"1810";
            when "01" & x"a6a" => DATA <= x"4f53";
            when "01" & x"a6b" => DATA <= x"5f43";
            when "01" & x"a6c" => DATA <= x"6f6e";
            when "01" & x"a6d" => DATA <= x"7665";
            when "01" & x"a6e" => DATA <= x"7274";
            when "01" & x"a6f" => DATA <= x"496e";
            when "01" & x"a70" => DATA <= x"7465";
            when "01" & x"a71" => DATA <= x"6765";
            when "01" & x"a72" => DATA <= x"7231";
            when "01" & x"a73" => DATA <= x"0000";
            when "01" & x"a74" => DATA <= x"0000";
            when "01" & x"a75" => DATA <= x"00da";
            when "01" & x"a76" => DATA <= x"003f";
            when "01" & x"a77" => DATA <= x"1838";
            when "01" & x"a78" => DATA <= x"4f53";
            when "01" & x"a79" => DATA <= x"5f43";
            when "01" & x"a7a" => DATA <= x"6f6e";
            when "01" & x"a7b" => DATA <= x"7665";
            when "01" & x"a7c" => DATA <= x"7274";
            when "01" & x"a7d" => DATA <= x"496e";
            when "01" & x"a7e" => DATA <= x"7465";
            when "01" & x"a7f" => DATA <= x"6765";
            when "01" & x"a80" => DATA <= x"7232";
            when "01" & x"a81" => DATA <= x"0000";
            when "01" & x"a82" => DATA <= x"0000";
            when "01" & x"a83" => DATA <= x"00db";
            when "01" & x"a84" => DATA <= x"003f";
            when "01" & x"a85" => DATA <= x"1860";
            when "01" & x"a86" => DATA <= x"4f53";
            when "01" & x"a87" => DATA <= x"5f43";
            when "01" & x"a88" => DATA <= x"6f6e";
            when "01" & x"a89" => DATA <= x"7665";
            when "01" & x"a8a" => DATA <= x"7274";
            when "01" & x"a8b" => DATA <= x"496e";
            when "01" & x"a8c" => DATA <= x"7465";
            when "01" & x"a8d" => DATA <= x"6765";
            when "01" & x"a8e" => DATA <= x"7233";
            when "01" & x"a8f" => DATA <= x"0000";
            when "01" & x"a90" => DATA <= x"0000";
            when "01" & x"a91" => DATA <= x"00dc";
            when "01" & x"a92" => DATA <= x"003f";
            when "01" & x"a93" => DATA <= x"1888";
            when "01" & x"a94" => DATA <= x"4f53";
            when "01" & x"a95" => DATA <= x"5f43";
            when "01" & x"a96" => DATA <= x"6f6e";
            when "01" & x"a97" => DATA <= x"7665";
            when "01" & x"a98" => DATA <= x"7274";
            when "01" & x"a99" => DATA <= x"496e";
            when "01" & x"a9a" => DATA <= x"7465";
            when "01" & x"a9b" => DATA <= x"6765";
            when "01" & x"a9c" => DATA <= x"7234";
            when "01" & x"a9d" => DATA <= x"0000";
            when "01" & x"a9e" => DATA <= x"0000";
            when "01" & x"a9f" => DATA <= x"00dd";
            when "01" & x"aa0" => DATA <= x"003f";
            when "01" & x"aa1" => DATA <= x"190a";
            when "01" & x"aa2" => DATA <= x"4f53";
            when "01" & x"aa3" => DATA <= x"5f43";
            when "01" & x"aa4" => DATA <= x"6f6e";
            when "01" & x"aa5" => DATA <= x"7665";
            when "01" & x"aa6" => DATA <= x"7274";
            when "01" & x"aa7" => DATA <= x"4269";
            when "01" & x"aa8" => DATA <= x"6e61";
            when "01" & x"aa9" => DATA <= x"7279";
            when "01" & x"aaa" => DATA <= x"3100";
            when "01" & x"aab" => DATA <= x"0000";
            when "01" & x"aac" => DATA <= x"0000";
            when "01" & x"aad" => DATA <= x"00de";
            when "01" & x"aae" => DATA <= x"003f";
            when "01" & x"aaf" => DATA <= x"1928";
            when "01" & x"ab0" => DATA <= x"4f53";
            when "01" & x"ab1" => DATA <= x"5f43";
            when "01" & x"ab2" => DATA <= x"6f6e";
            when "01" & x"ab3" => DATA <= x"7665";
            when "01" & x"ab4" => DATA <= x"7274";
            when "01" & x"ab5" => DATA <= x"4269";
            when "01" & x"ab6" => DATA <= x"6e61";
            when "01" & x"ab7" => DATA <= x"7279";
            when "01" & x"ab8" => DATA <= x"3200";
            when "01" & x"ab9" => DATA <= x"0000";
            when "01" & x"aba" => DATA <= x"0000";
            when "01" & x"abb" => DATA <= x"00df";
            when "01" & x"abc" => DATA <= x"003f";
            when "01" & x"abd" => DATA <= x"1948";
            when "01" & x"abe" => DATA <= x"4f53";
            when "01" & x"abf" => DATA <= x"5f43";
            when "01" & x"ac0" => DATA <= x"6f6e";
            when "01" & x"ac1" => DATA <= x"7665";
            when "01" & x"ac2" => DATA <= x"7274";
            when "01" & x"ac3" => DATA <= x"4269";
            when "01" & x"ac4" => DATA <= x"6e61";
            when "01" & x"ac5" => DATA <= x"7279";
            when "01" & x"ac6" => DATA <= x"3300";
            when "01" & x"ac7" => DATA <= x"0000";
            when "01" & x"ac8" => DATA <= x"0000";
            when "01" & x"ac9" => DATA <= x"00e0";
            when "01" & x"aca" => DATA <= x"003f";
            when "01" & x"acb" => DATA <= x"1966";
            when "01" & x"acc" => DATA <= x"4f53";
            when "01" & x"acd" => DATA <= x"5f43";
            when "01" & x"ace" => DATA <= x"6f6e";
            when "01" & x"acf" => DATA <= x"7665";
            when "01" & x"ad0" => DATA <= x"7274";
            when "01" & x"ad1" => DATA <= x"4269";
            when "01" & x"ad2" => DATA <= x"6e61";
            when "01" & x"ad3" => DATA <= x"7279";
            when "01" & x"ad4" => DATA <= x"3400";
            when "01" & x"ad5" => DATA <= x"0000";
            when "01" & x"ad6" => DATA <= x"0000";
            when "01" & x"ad7" => DATA <= x"00ea";
            when "01" & x"ad8" => DATA <= x"003f";
            when "01" & x"ad9" => DATA <= x"19e2";
            when "01" & x"ada" => DATA <= x"4f53";
            when "01" & x"adb" => DATA <= x"5f43";
            when "01" & x"adc" => DATA <= x"6f6e";
            when "01" & x"add" => DATA <= x"7665";
            when "01" & x"ade" => DATA <= x"7274";
            when "01" & x"adf" => DATA <= x"4e65";
            when "01" & x"ae0" => DATA <= x"7453";
            when "01" & x"ae1" => DATA <= x"7461";
            when "01" & x"ae2" => DATA <= x"7469";
            when "01" & x"ae3" => DATA <= x"6f6e";
            when "01" & x"ae4" => DATA <= x"0000";
            when "01" & x"ae5" => DATA <= x"00ff";
            when "01" & x"ae6" => DATA <= x"003f";
            when "01" & x"ae7" => DATA <= x"1b52";
            when "01" & x"ae8" => DATA <= x"4552";
            when "01" & x"ae9" => DATA <= x"524f";
            when "01" & x"aea" => DATA <= x"5220";
            when "01" & x"aeb" => DATA <= x"2000";
            when "01" & x"aec" => DATA <= x"003f";
            when "01" & x"aed" => DATA <= x"1bb0";
            when "01" & x"aee" => DATA <= x"464c";
            when "01" & x"aef" => DATA <= x"4153";
            when "01" & x"af0" => DATA <= x"4820";
            when "01" & x"af1" => DATA <= x"2000";
            when "01" & x"af2" => DATA <= x"003f";
            when "01" & x"af3" => DATA <= x"1c88";
            when "01" & x"af4" => DATA <= x"474f";
            when "01" & x"af5" => DATA <= x"2000";
            when "01" & x"af6" => DATA <= x"003f";
            when "01" & x"af7" => DATA <= x"1cb6";
            when "01" & x"af8" => DATA <= x"4845";
            when "01" & x"af9" => DATA <= x"4c50";
            when "01" & x"afa" => DATA <= x"2020";
            when "01" & x"afb" => DATA <= x"2000";
            when "01" & x"afc" => DATA <= x"003f";
            when "01" & x"afd" => DATA <= x"1db2";
            when "01" & x"afe" => DATA <= x"4d4f";
            when "01" & x"aff" => DATA <= x"4e00";
            when "01" & x"b00" => DATA <= x"003f";
            when "01" & x"b01" => DATA <= x"247c";
            when "01" & x"b02" => DATA <= x"5155";
            when "01" & x"b03" => DATA <= x"4954";
            when "01" & x"b04" => DATA <= x"2020";
            when "01" & x"b05" => DATA <= x"2000";
            when "01" & x"b06" => DATA <= x"003f";
            when "01" & x"b07" => DATA <= x"2480";
            when "01" & x"b08" => DATA <= x"545a";
            when "01" & x"b09" => DATA <= x"4150";
            when "01" & x"b0a" => DATA <= x"2020";
            when "01" & x"b0b" => DATA <= x"2000";
            when "01" & x"b0c" => DATA <= x"003f";
            when "01" & x"b0d" => DATA <= x"2484";
            when "01" & x"b0e" => DATA <= x"5846";
            when "01" & x"b0f" => DATA <= x"4552";
            when "01" & x"b10" => DATA <= x"2020";
            when "01" & x"b11" => DATA <= x"2000";
            when "01" & x"b12" => DATA <= x"ffff";
            when "01" & x"b13" => DATA <= x"ffff";
            when "01" & x"b14" => DATA <= x"0000";
            when "01" & x"b15" => DATA <= x"0508";
            when "01" & x"b16" => DATA <= x"0000";
            when "01" & x"b17" => DATA <= x"0508";
            when "01" & x"b18" => DATA <= x"0000";
            when "01" & x"b19" => DATA <= x"0000";
            when "01" & x"b1a" => DATA <= x"0000";
            when "01" & x"b1b" => DATA <= x"0000";
            when "01" & x"b1c" => DATA <= x"0000";
            when "01" & x"b1d" => DATA <= x"0010";
            when "01" & x"b1e" => DATA <= x"0000";
            when "01" & x"b1f" => DATA <= x"0000";
            when "01" & x"b20" => DATA <= x"0000";
            when "01" & x"b21" => DATA <= x"0000";
            when "01" & x"b22" => DATA <= x"0000";
            when "01" & x"b23" => DATA <= x"0000";
            when "01" & x"b24" => DATA <= x"0000";
            when "01" & x"b25" => DATA <= x"0000";
            when "01" & x"b26" => DATA <= x"0000";
            when "01" & x"b27" => DATA <= x"0000";
            when "01" & x"b28" => DATA <= x"0000";
            when "01" & x"b29" => DATA <= x"0000";
            when "01" & x"b2a" => DATA <= x"0000";
            when "01" & x"b2b" => DATA <= x"0000";
            when "01" & x"b2c" => DATA <= x"0000";
            when "01" & x"b2d" => DATA <= x"0000";
            when "01" & x"b2e" => DATA <= x"0000";
            when "01" & x"b2f" => DATA <= x"000c";
            when "01" & x"b30" => DATA <= x"0000";
            when "01" & x"b31" => DATA <= x"0000";
            when "01" & x"b32" => DATA <= x"0000";
            when "01" & x"b33" => DATA <= x"0000";
            when "01" & x"b34" => DATA <= x"0000";
            when "01" & x"b35" => DATA <= x"04c0";
            when "01" & x"b36" => DATA <= x"0000";
            when "01" & x"b37" => DATA <= x"0000";
            when "01" & x"b38" => DATA <= x"0000";
            when "01" & x"b39" => DATA <= x"0000";
            when "01" & x"b3a" => DATA <= x"0000";
            when "01" & x"b3b" => DATA <= x"0404";
            when "01" & x"b3c" => DATA <= x"0000";
            when "01" & x"b3d" => DATA <= x"04d4";
            when "01" & x"b3e" => DATA <= x"0000";
            when "01" & x"b3f" => DATA <= x"04f4";
            when "01" & x"b40" => DATA <= x"0000";
            when "01" & x"b41" => DATA <= x"04c4";
            when "01" & x"b42" => DATA <= x"0000";
            when "01" & x"b43" => DATA <= x"04d8";
            when "01" & x"b44" => DATA <= x"0000";
            when "01" & x"b45" => DATA <= x"04f8";
            when "01" & x"b46" => DATA <= x"0000";
            when "01" & x"b47" => DATA <= x"04c8";
            when "01" & x"b48" => DATA <= x"0000";
            when "01" & x"b49" => DATA <= x"04dc";
            when "01" & x"b4a" => DATA <= x"0000";
            when "01" & x"b4b" => DATA <= x"04fc";
            when "01" & x"b4c" => DATA <= x"0000";
            when "01" & x"b4d" => DATA <= x"04cc";
            when "01" & x"b4e" => DATA <= x"0000";
            when "01" & x"b4f" => DATA <= x"04e0";
            when "01" & x"b50" => DATA <= x"0000";
            when "01" & x"b51" => DATA <= x"0000";
            when "01" & x"b52" => DATA <= x"0000";
            when "01" & x"b53" => DATA <= x"0440";
            when "01" & x"b54" => DATA <= x"0000";
            when "01" & x"b55" => DATA <= x"04e4";
            when "01" & x"b56" => DATA <= x"0000";
            when "01" & x"b57" => DATA <= x"0000";
            when "01" & x"b58" => DATA <= x"0000";
            when "01" & x"b59" => DATA <= x"04d0";
            when "01" & x"b5a" => DATA <= x"0000";
            when "01" & x"b5b" => DATA <= x"04e8";
            when "01" & x"b5c" => DATA <= x"0000";
            when "01" & x"b5d" => DATA <= x"0000";
            when "01" & x"b5e" => DATA <= x"0000";
            when "01" & x"b5f" => DATA <= x"0460";
            when "01" & x"b60" => DATA <= x"0000";
            when "01" & x"b61" => DATA <= x"04ec";
            when "01" & x"b62" => DATA <= x"0000";
            when "01" & x"b63" => DATA <= x"0000";
            when "01" & x"b64" => DATA <= x"0000";
            when "01" & x"b65" => DATA <= x"0538";
            when "01" & x"b66" => DATA <= x"0000";
            when "01" & x"b67" => DATA <= x"0000";
            when "01" & x"b68" => DATA <= x"0000";
            when "01" & x"b69" => DATA <= x"0000";
            when "01" & x"b6a" => DATA <= x"0000";
            when "01" & x"b6b" => DATA <= x"050c";
            when "01" & x"b6c" => DATA <= x"0000";
            when "01" & x"b6d" => DATA <= x"0000";
            when "01" & x"b6e" => DATA <= x"0000";
            when "01" & x"b6f" => DATA <= x"0000";
            when "01" & x"b70" => DATA <= x"0000";
            when "01" & x"b71" => DATA <= x"0000";
            when "01" & x"b72" => DATA <= x"0000";
            when "01" & x"b73" => DATA <= x"0000";
            when "01" & x"b74" => DATA <= x"0000";
            when "01" & x"b75" => DATA <= x"0000";
            when "01" & x"b76" => DATA <= x"0000";
            when "01" & x"b77" => DATA <= x"0474";
            when "01" & x"b78" => DATA <= x"0000";
            when "01" & x"b79" => DATA <= x"04f0";
            when "01" & x"b7a" => DATA <= x"0000";
            when "01" & x"b7b" => DATA <= x"0000";
            when "01" & x"b7c" => DATA <= x"003f";
            when "01" & x"b7d" => DATA <= x"0776";
            when "01" & x"b7e" => DATA <= x"003f";
            when "01" & x"b7f" => DATA <= x"0776";
            when "01" & x"b80" => DATA <= x"003f";
            when "01" & x"b81" => DATA <= x"0776";
            when "01" & x"b82" => DATA <= x"003f";
            when "01" & x"b83" => DATA <= x"0776";
            when "01" & x"b84" => DATA <= x"003f";
            when "01" & x"b85" => DATA <= x"0776";
            when "01" & x"b86" => DATA <= x"003f";
            when "01" & x"b87" => DATA <= x"0776";
            when "01" & x"b88" => DATA <= x"003f";
            when "01" & x"b89" => DATA <= x"0776";
            when "01" & x"b8a" => DATA <= x"003f";
            when "01" & x"b8b" => DATA <= x"0776";
            when "01" & x"b8c" => DATA <= x"003f";
            when "01" & x"b8d" => DATA <= x"0776";
            when "01" & x"b8e" => DATA <= x"003f";
            when "01" & x"b8f" => DATA <= x"0776";
            when "01" & x"b90" => DATA <= x"003f";
            when "01" & x"b91" => DATA <= x"1104";
            when "01" & x"b92" => DATA <= x"003f";
            when "01" & x"b93" => DATA <= x"0776";
            when "01" & x"b94" => DATA <= x"003f";
            when "01" & x"b95" => DATA <= x"0776";
            when "01" & x"b96" => DATA <= x"003f";
            when "01" & x"b97" => DATA <= x"0776";
            when "01" & x"b98" => DATA <= x"003f";
            when "01" & x"b99" => DATA <= x"0776";
            when "01" & x"b9a" => DATA <= x"003f";
            when "01" & x"b9b" => DATA <= x"0776";
            when "01" & x"b9c" => DATA <= x"003f";
            when "01" & x"b9d" => DATA <= x"0776";
            when "01" & x"b9e" => DATA <= x"003f";
            when "01" & x"b9f" => DATA <= x"0776";
            when "01" & x"ba0" => DATA <= x"003f";
            when "01" & x"ba1" => DATA <= x"0776";
            when "01" & x"ba2" => DATA <= x"003f";
            when "01" & x"ba3" => DATA <= x"0776";
            when "01" & x"ba4" => DATA <= x"003f";
            when "01" & x"ba5" => DATA <= x"0776";
            when "01" & x"ba6" => DATA <= x"003f";
            when "01" & x"ba7" => DATA <= x"0776";
            when "01" & x"ba8" => DATA <= x"003f";
            when "01" & x"ba9" => DATA <= x"1112";
            when "01" & x"baa" => DATA <= x"003f";
            when "01" & x"bab" => DATA <= x"0776";
            when "01" & x"bac" => DATA <= x"003f";
            when "01" & x"bad" => DATA <= x"0776";
            when "01" & x"bae" => DATA <= x"003f";
            when "01" & x"baf" => DATA <= x"0776";
            when "01" & x"bb0" => DATA <= x"003f";
            when "01" & x"bb1" => DATA <= x"0776";
            when "01" & x"bb2" => DATA <= x"003f";
            when "01" & x"bb3" => DATA <= x"0776";
            when "01" & x"bb4" => DATA <= x"003f";
            when "01" & x"bb5" => DATA <= x"0776";
            when "01" & x"bb6" => DATA <= x"003f";
            when "01" & x"bb7" => DATA <= x"0776";
            when "01" & x"bb8" => DATA <= x"003f";
            when "01" & x"bb9" => DATA <= x"0776";
            when "01" & x"bba" => DATA <= x"003f";
            when "01" & x"bbb" => DATA <= x"0776";
            when "01" & x"bbc" => DATA <= x"003f";
            when "01" & x"bbd" => DATA <= x"0776";
            when "01" & x"bbe" => DATA <= x"003f";
            when "01" & x"bbf" => DATA <= x"0776";
            when "01" & x"bc0" => DATA <= x"003f";
            when "01" & x"bc1" => DATA <= x"0776";
            when "01" & x"bc2" => DATA <= x"003f";
            when "01" & x"bc3" => DATA <= x"0776";
            when "01" & x"bc4" => DATA <= x"003f";
            when "01" & x"bc5" => DATA <= x"0776";
            when "01" & x"bc6" => DATA <= x"003f";
            when "01" & x"bc7" => DATA <= x"0776";
            when "01" & x"bc8" => DATA <= x"003f";
            when "01" & x"bc9" => DATA <= x"0776";
            when "01" & x"bca" => DATA <= x"003f";
            when "01" & x"bcb" => DATA <= x"0776";
            when "01" & x"bcc" => DATA <= x"003f";
            when "01" & x"bcd" => DATA <= x"0776";
            when "01" & x"bce" => DATA <= x"003f";
            when "01" & x"bcf" => DATA <= x"0776";
            when "01" & x"bd0" => DATA <= x"003f";
            when "01" & x"bd1" => DATA <= x"0776";
            when "01" & x"bd2" => DATA <= x"003f";
            when "01" & x"bd3" => DATA <= x"0776";
            when "01" & x"bd4" => DATA <= x"003f";
            when "01" & x"bd5" => DATA <= x"0776";
            when "01" & x"bd6" => DATA <= x"003f";
            when "01" & x"bd7" => DATA <= x"0776";
            when "01" & x"bd8" => DATA <= x"003f";
            when "01" & x"bd9" => DATA <= x"0776";
            when "01" & x"bda" => DATA <= x"003f";
            when "01" & x"bdb" => DATA <= x"0776";
            when "01" & x"bdc" => DATA <= x"003f";
            when "01" & x"bdd" => DATA <= x"0776";
            when "01" & x"bde" => DATA <= x"003f";
            when "01" & x"bdf" => DATA <= x"0776";
            when "01" & x"be0" => DATA <= x"003f";
            when "01" & x"be1" => DATA <= x"0776";
            when "01" & x"be2" => DATA <= x"003f";
            when "01" & x"be3" => DATA <= x"0776";
            when "01" & x"be4" => DATA <= x"003f";
            when "01" & x"be5" => DATA <= x"0776";
            when "01" & x"be6" => DATA <= x"003f";
            when "01" & x"be7" => DATA <= x"0776";
            when "01" & x"be8" => DATA <= x"003f";
            when "01" & x"be9" => DATA <= x"0776";
            when "01" & x"bea" => DATA <= x"003f";
            when "01" & x"beb" => DATA <= x"0776";
            when "01" & x"bec" => DATA <= x"003f";
            when "01" & x"bed" => DATA <= x"0776";
            when "01" & x"bee" => DATA <= x"003f";
            when "01" & x"bef" => DATA <= x"0776";
            when "01" & x"bf0" => DATA <= x"003f";
            when "01" & x"bf1" => DATA <= x"0776";
            when "01" & x"bf2" => DATA <= x"1890";
            when "01" & x"bf3" => DATA <= x"0210";
            when "01" & x"bf4" => DATA <= x"e3c9";
            when "01" & x"bf5" => DATA <= x"faf0";
            when "01" & x"bf6" => DATA <= x"036c";
            when "01" & x"bf7" => DATA <= x"0325";
            when "01" & x"bf8" => DATA <= x"8670";
            when "01" & x"bf9" => DATA <= x"8471";
            when "01" & x"bfa" => DATA <= x"48a9";
            when "01" & x"bfb" => DATA <= x"fba2";
            when "01" & x"bfc" => DATA <= x"00a0";
            when "01" & x"bfd" => DATA <= x"ff20";
            when "01" & x"bfe" => DATA <= x"f4ff";
            when "01" & x"bff" => DATA <= x"8673";
            when "01" & x"c00" => DATA <= x"ad34";
            when "01" & x"c01" => DATA <= x"fe48";
            when "01" & x"c02" => DATA <= x"a9c7";
            when "01" & x"c03" => DATA <= x"2006";
            when "01" & x"c04" => DATA <= x"0490";
            when "01" & x"c05" => DATA <= x"f9a0";
            when "01" & x"c06" => DATA <= x"00b1";
            when "01" & x"c07" => DATA <= x"70c9";
            when "01" & x"c08" => DATA <= x"0d08";
            when "01" & x"c09" => DATA <= x"a5f4";
            when "01" & x"c0a" => DATA <= x"8572";
            when "01" & x"c0b" => DATA <= x"a00d";
            when "01" & x"c0c" => DATA <= x"b170";
            when "01" & x"c0d" => DATA <= x"aaa0";
            when "01" & x"c0e" => DATA <= x"02b1";
            when "01" & x"c0f" => DATA <= x"7085";
            when "01" & x"c10" => DATA <= x"74c8";
            when "01" & x"c11" => DATA <= x"b170";
            when "01" & x"c12" => DATA <= x"8575";
            when "01" & x"c13" => DATA <= x"28f0";
            when "01" & x"c14" => DATA <= x"408a";
            when "01" & x"c15" => DATA <= x"4829";
            when "01" & x"c16" => DATA <= x"40d0";
            when "01" & x"c17" => DATA <= x"138a";
            when "01" & x"c18" => DATA <= x"2920";
            when "01" & x"c19" => DATA <= x"d004";
            when "01" & x"c1a" => DATA <= x"a200";
            when "01" & x"c1b" => DATA <= x"f002";
            when "01" & x"c1c" => DATA <= x"a201";
            when "01" & x"c1d" => DATA <= x"a96c";
            when "01" & x"c1e" => DATA <= x"20f4";
            when "01" & x"c1f" => DATA <= x"ff4c";
            when "01" & x"c20" => DATA <= x"7725";
            when "01" & x"c21" => DATA <= x"a984";
            when "01" & x"c22" => DATA <= x"20f4";
            when "01" & x"c23" => DATA <= x"ffc0";
            when "01" & x"c24" => DATA <= x"80d0";
            when "01" & x"c25" => DATA <= x"08a9";
            when "01" & x"c26" => DATA <= x"01c5";
            when "01" & x"c27" => DATA <= x"73d0";
            when "01" & x"c28" => DATA <= x"e7f0";
            when "01" & x"c29" => DATA <= x"e1a9";
            when "01" & x"c2a" => DATA <= x"02c5";
            when "01" & x"c2b" => DATA <= x"73d0";
            when "01" & x"c2c" => DATA <= x"dbf0";
            when "01" & x"c2d" => DATA <= x"dd68";
            when "01" & x"c2e" => DATA <= x"aa29";
            when "01" & x"c2f" => DATA <= x"10d0";
            when "01" & x"c30" => DATA <= x"088a";
            when "01" & x"c31" => DATA <= x"290f";
            when "01" & x"c32" => DATA <= x"85f4";
            when "01" & x"c33" => DATA <= x"8d30";
            when "01" & x"c34" => DATA <= x"fea0";
            when "01" & x"c35" => DATA <= x"0ab1";
            when "01" & x"c36" => DATA <= x"7085";
            when "01" & x"c37" => DATA <= x"77c8";
            when "01" & x"c38" => DATA <= x"b170";
            when "01" & x"c39" => DATA <= x"8576";
            when "01" & x"c3a" => DATA <= x"0577";
            when "01" & x"c3b" => DATA <= x"d002";
            when "01" & x"c3c" => DATA <= x"f06e";
            when "01" & x"c3d" => DATA <= x"a577";
            when "01" & x"c3e" => DATA <= x"f002";
            when "01" & x"c3f" => DATA <= x"e676";
            when "01" & x"c40" => DATA <= x"c8b1";
            when "01" & x"c41" => DATA <= x"7048";
            when "01" & x"c42" => DATA <= x"a577";
            when "01" & x"c43" => DATA <= x"f011";
            when "01" & x"c44" => DATA <= x"a576";
            when "01" & x"c45" => DATA <= x"c901";
            when "01" & x"c46" => DATA <= x"d00b";
            when "01" & x"c47" => DATA <= x"6848";
            when "01" & x"c48" => DATA <= x"c906";
            when "01" & x"c49" => DATA <= x"9005";
            when "01" & x"c4a" => DATA <= x"6838";
            when "01" & x"c4b" => DATA <= x"e906";
            when "01" & x"c4c" => DATA <= x"48a5";
            when "01" & x"c4d" => DATA <= x"7018";
            when "01" & x"c4e" => DATA <= x"6906";
            when "01" & x"c4f" => DATA <= x"aaa9";
            when "01" & x"c50" => DATA <= x"0065";
            when "01" & x"c51" => DATA <= x"71a8";
            when "01" & x"c52" => DATA <= x"6848";
            when "01" & x"c53" => DATA <= x"2006";
            when "01" & x"c54" => DATA <= x"04a6";
            when "01" & x"c55" => DATA <= x"7768";
            when "01" & x"c56" => DATA <= x"a000";
            when "01" & x"c57" => DATA <= x"c900";
            when "01" & x"c58" => DATA <= x"f01e";
            when "01" & x"c59" => DATA <= x"c901";
            when "01" & x"c5a" => DATA <= x"f035";
            when "01" & x"c5b" => DATA <= x"c902";
            when "01" & x"c5c" => DATA <= x"f049";
            when "01" & x"c5d" => DATA <= x"c903";
            when "01" & x"c5e" => DATA <= x"f070";
            when "01" & x"c5f" => DATA <= x"c906";
            when "01" & x"c60" => DATA <= x"f008";
            when "01" & x"c61" => DATA <= x"c907";
            when "01" & x"c62" => DATA <= x"f007";
            when "01" & x"c63" => DATA <= x"a900";
            when "01" & x"c64" => DATA <= x"f01e";
            when "01" & x"c65" => DATA <= x"4c75";
            when "01" & x"c66" => DATA <= x"264c";
            when "01" & x"c67" => DATA <= x"a326";
            when "01" & x"c68" => DATA <= x"20f4";
            when "01" & x"c69" => DATA <= x"26ad";
            when "01" & x"c6a" => DATA <= x"e5fe";
            when "01" & x"c6b" => DATA <= x"9174";
            when "01" & x"c6c" => DATA <= x"20f4";
            when "01" & x"c6d" => DATA <= x"26e6";
            when "01" & x"c6e" => DATA <= x"74d0";
            when "01" & x"c6f" => DATA <= x"02e6";
            when "01" & x"c70" => DATA <= x"75ca";
            when "01" & x"c71" => DATA <= x"d0ef";
            when "01" & x"c72" => DATA <= x"c676";
            when "01" & x"c73" => DATA <= x"d0eb";
            when "01" & x"c74" => DATA <= x"4cda";
            when "01" & x"c75" => DATA <= x"26b1";
            when "01" & x"c76" => DATA <= x"748d";
            when "01" & x"c77" => DATA <= x"e5fe";
            when "01" & x"c78" => DATA <= x"20f4";
            when "01" & x"c79" => DATA <= x"26e6";
            when "01" & x"c7a" => DATA <= x"74d0";
            when "01" & x"c7b" => DATA <= x"02e6";
            when "01" & x"c7c" => DATA <= x"75ca";
            when "01" & x"c7d" => DATA <= x"d0ef";
            when "01" & x"c7e" => DATA <= x"c676";
            when "01" & x"c7f" => DATA <= x"d0eb";
            when "01" & x"c80" => DATA <= x"4cda";
            when "01" & x"c81" => DATA <= x"2620";
            when "01" & x"c82" => DATA <= x"f426";
            when "01" & x"c83" => DATA <= x"ade5";
            when "01" & x"c84" => DATA <= x"fe91";
            when "01" & x"c85" => DATA <= x"74e6";
            when "01" & x"c86" => DATA <= x"74d0";
            when "01" & x"c87" => DATA <= x"02e6";
            when "01" & x"c88" => DATA <= x"75ea";
            when "01" & x"c89" => DATA <= x"eaad";
            when "01" & x"c8a" => DATA <= x"e5fe";
            when "01" & x"c8b" => DATA <= x"9174";
            when "01" & x"c8c" => DATA <= x"e674";
            when "01" & x"c8d" => DATA <= x"d002";
            when "01" & x"c8e" => DATA <= x"e675";
            when "01" & x"c8f" => DATA <= x"20f3";
            when "01" & x"c90" => DATA <= x"26ea";
            when "01" & x"c91" => DATA <= x"eaca";
            when "01" & x"c92" => DATA <= x"cad0";
            when "01" & x"c93" => DATA <= x"dfc6";
            when "01" & x"c94" => DATA <= x"76d0";
            when "01" & x"c95" => DATA <= x"db4c";
            when "01" & x"c96" => DATA <= x"da26";
            when "01" & x"c97" => DATA <= x"b174";
            when "01" & x"c98" => DATA <= x"8de5";
            when "01" & x"c99" => DATA <= x"fee6";
            when "01" & x"c9a" => DATA <= x"74f0";
            when "01" & x"c9b" => DATA <= x"03ea";
            when "01" & x"c9c" => DATA <= x"d002";
            when "01" & x"c9d" => DATA <= x"e675";
            when "01" & x"c9e" => DATA <= x"a573";
            when "01" & x"c9f" => DATA <= x"b174";
            when "01" & x"ca0" => DATA <= x"8de5";
            when "01" & x"ca1" => DATA <= x"fee6";
            when "01" & x"ca2" => DATA <= x"74f0";
            when "01" & x"ca3" => DATA <= x"03ea";
            when "01" & x"ca4" => DATA <= x"d002";
            when "01" & x"ca5" => DATA <= x"e675";
            when "01" & x"ca6" => DATA <= x"20f3";
            when "01" & x"ca7" => DATA <= x"26ca";
            when "01" & x"ca8" => DATA <= x"cad0";
            when "01" & x"ca9" => DATA <= x"dbc6";
            when "01" & x"caa" => DATA <= x"76d0";
            when "01" & x"cab" => DATA <= x"d7f0";
            when "01" & x"cac" => DATA <= x"6520";
            when "01" & x"cad" => DATA <= x"f426";
            when "01" & x"cae" => DATA <= x"ade5";
            when "01" & x"caf" => DATA <= x"fe91";
            when "01" & x"cb0" => DATA <= x"74ea";
            when "01" & x"cb1" => DATA <= x"eaea";
            when "01" & x"cb2" => DATA <= x"c8d0";
            when "01" & x"cb3" => DATA <= x"f5e0";
            when "01" & x"cb4" => DATA <= x"00d0";
            when "01" & x"cb5" => DATA <= x"0cc6";
            when "01" & x"cb6" => DATA <= x"76f0";
            when "01" & x"cb7" => DATA <= x"4f20";
            when "01" & x"cb8" => DATA <= x"ce26";
            when "01" & x"cb9" => DATA <= x"a906";
            when "01" & x"cba" => DATA <= x"4c9f";
            when "01" & x"cbb" => DATA <= x"25c6";
            when "01" & x"cbc" => DATA <= x"76a5";
            when "01" & x"cbd" => DATA <= x"76c9";
            when "01" & x"cbe" => DATA <= x"01d0";
            when "01" & x"cbf" => DATA <= x"f020";
            when "01" & x"cc0" => DATA <= x"ce26";
            when "01" & x"cc1" => DATA <= x"a900";
            when "01" & x"cc2" => DATA <= x"4c9f";
            when "01" & x"cc3" => DATA <= x"25b1";
            when "01" & x"cc4" => DATA <= x"748d";
            when "01" & x"cc5" => DATA <= x"e5fe";
            when "01" & x"cc6" => DATA <= x"eaea";
            when "01" & x"cc7" => DATA <= x"eac8";
            when "01" & x"cc8" => DATA <= x"d0f5";
            when "01" & x"cc9" => DATA <= x"e000";
            when "01" & x"cca" => DATA <= x"d00c";
            when "01" & x"ccb" => DATA <= x"c676";
            when "01" & x"ccc" => DATA <= x"f024";
            when "01" & x"ccd" => DATA <= x"20ce";
            when "01" & x"cce" => DATA <= x"26a9";
            when "01" & x"ccf" => DATA <= x"074c";
            when "01" & x"cd0" => DATA <= x"9f25";
            when "01" & x"cd1" => DATA <= x"c676";
            when "01" & x"cd2" => DATA <= x"a576";
            when "01" & x"cd3" => DATA <= x"c901";
            when "01" & x"cd4" => DATA <= x"d0f0";
            when "01" & x"cd5" => DATA <= x"20ce";
            when "01" & x"cd6" => DATA <= x"26a9";
            when "01" & x"cd7" => DATA <= x"014c";
            when "01" & x"cd8" => DATA <= x"9f25";
            when "01" & x"cd9" => DATA <= x"e675";
            when "01" & x"cda" => DATA <= x"a007";
            when "01" & x"cdb" => DATA <= x"b170";
            when "01" & x"cdc" => DATA <= x"1869";
            when "01" & x"cdd" => DATA <= x"0191";
            when "01" & x"cde" => DATA <= x"7060";
            when "01" & x"cdf" => DATA <= x"a987";
            when "01" & x"ce0" => DATA <= x"2006";
            when "01" & x"ce1" => DATA <= x"04a5";
            when "01" & x"ce2" => DATA <= x"72c5";
            when "01" & x"ce3" => DATA <= x"f4f0";
            when "01" & x"ce4" => DATA <= x"0585";
            when "01" & x"ce5" => DATA <= x"f48d";
            when "01" & x"ce6" => DATA <= x"30fe";
            when "01" & x"ce7" => DATA <= x"688d";
            when "01" & x"ce8" => DATA <= x"34fe";
            when "01" & x"ce9" => DATA <= x"a670";
            when "01" & x"cea" => DATA <= x"a471";
            when "01" & x"ceb" => DATA <= x"6860";
            when "01" & x"cec" => DATA <= x"20f3";
            when "01" & x"ced" => DATA <= x"2620";
            when "01" & x"cee" => DATA <= x"f326";
            when "01" & x"cef" => DATA <= x"60ff";
            when "01" & x"cf0" => DATA <= x"003c";
            when "01" & x"cf1" => DATA <= x"ffff";
            when "01" & x"cf2" => DATA <= x"4f52";
            when "01" & x"cf3" => DATA <= x"4920";
            when "01" & x"cf4" => DATA <= x"2000";
            when "01" & x"cf5" => DATA <= x"003f";
            when "01" & x"cf6" => DATA <= x"39e0";
            when "01" & x"cf7" => DATA <= x"007c";
            when "01" & x"cf8" => DATA <= x"ffff";
            when "01" & x"cf9" => DATA <= x"4f52";
            when "01" & x"cfa" => DATA <= x"4920";
            when "01" & x"cfb" => DATA <= x"2000";
            when "01" & x"cfc" => DATA <= x"003f";
            when "01" & x"cfd" => DATA <= x"39e0";
            when "01" & x"cfe" => DATA <= x"023c";
            when "01" & x"cff" => DATA <= x"ffff";
            when "01" & x"d00" => DATA <= x"414e";
            when "01" & x"d01" => DATA <= x"4449";
            when "01" & x"d02" => DATA <= x"2000";
            when "01" & x"d03" => DATA <= x"003f";
            when "01" & x"d04" => DATA <= x"39e0";
            when "01" & x"d05" => DATA <= x"027c";
            when "01" & x"d06" => DATA <= x"ffff";
            when "01" & x"d07" => DATA <= x"414e";
            when "01" & x"d08" => DATA <= x"4449";
            when "01" & x"d09" => DATA <= x"2000";
            when "01" & x"d0a" => DATA <= x"003f";
            when "01" & x"d0b" => DATA <= x"39e0";
            when "01" & x"d0c" => DATA <= x"0a3c";
            when "01" & x"d0d" => DATA <= x"ffff";
            when "01" & x"d0e" => DATA <= x"454f";
            when "01" & x"d0f" => DATA <= x"5249";
            when "01" & x"d10" => DATA <= x"2000";
            when "01" & x"d11" => DATA <= x"003f";
            when "01" & x"d12" => DATA <= x"39e0";
            when "01" & x"d13" => DATA <= x"0a7c";
            when "01" & x"d14" => DATA <= x"ffff";
            when "01" & x"d15" => DATA <= x"454f";
            when "01" & x"d16" => DATA <= x"5249";
            when "01" & x"d17" => DATA <= x"2000";
            when "01" & x"d18" => DATA <= x"003f";
            when "01" & x"d19" => DATA <= x"39e0";
            when "01" & x"d1a" => DATA <= x"0800";
            when "01" & x"d1b" => DATA <= x"ffc0";
            when "01" & x"d1c" => DATA <= x"4254";
            when "01" & x"d1d" => DATA <= x"5354";
            when "01" & x"d1e" => DATA <= x"2000";
            when "01" & x"d1f" => DATA <= x"003f";
            when "01" & x"d20" => DATA <= x"39e0";
            when "01" & x"d21" => DATA <= x"0840";
            when "01" & x"d22" => DATA <= x"ffc0";
            when "01" & x"d23" => DATA <= x"4243";
            when "01" & x"d24" => DATA <= x"4847";
            when "01" & x"d25" => DATA <= x"2000";
            when "01" & x"d26" => DATA <= x"003f";
            when "01" & x"d27" => DATA <= x"39e0";
            when "01" & x"d28" => DATA <= x"0880";
            when "01" & x"d29" => DATA <= x"ffc0";
            when "01" & x"d2a" => DATA <= x"4243";
            when "01" & x"d2b" => DATA <= x"4c52";
            when "01" & x"d2c" => DATA <= x"2000";
            when "01" & x"d2d" => DATA <= x"003f";
            when "01" & x"d2e" => DATA <= x"39e0";
            when "01" & x"d2f" => DATA <= x"08c0";
            when "01" & x"d30" => DATA <= x"ffc0";
            when "01" & x"d31" => DATA <= x"4253";
            when "01" & x"d32" => DATA <= x"4554";
            when "01" & x"d33" => DATA <= x"2000";
            when "01" & x"d34" => DATA <= x"003f";
            when "01" & x"d35" => DATA <= x"39e0";
            when "01" & x"d36" => DATA <= x"0000";
            when "01" & x"d37" => DATA <= x"ff00";
            when "01" & x"d38" => DATA <= x"4f52";
            when "01" & x"d39" => DATA <= x"4920";
            when "01" & x"d3a" => DATA <= x"2000";
            when "01" & x"d3b" => DATA <= x"003f";
            when "01" & x"d3c" => DATA <= x"39e0";
            when "01" & x"d3d" => DATA <= x"0200";
            when "01" & x"d3e" => DATA <= x"ff00";
            when "01" & x"d3f" => DATA <= x"414e";
            when "01" & x"d40" => DATA <= x"4449";
            when "01" & x"d41" => DATA <= x"2000";
            when "01" & x"d42" => DATA <= x"003f";
            when "01" & x"d43" => DATA <= x"39e0";
            when "01" & x"d44" => DATA <= x"0400";
            when "01" & x"d45" => DATA <= x"ff00";
            when "01" & x"d46" => DATA <= x"5355";
            when "01" & x"d47" => DATA <= x"4249";
            when "01" & x"d48" => DATA <= x"2000";
            when "01" & x"d49" => DATA <= x"003f";
            when "01" & x"d4a" => DATA <= x"39e0";
            when "01" & x"d4b" => DATA <= x"0600";
            when "01" & x"d4c" => DATA <= x"ff00";
            when "01" & x"d4d" => DATA <= x"4144";
            when "01" & x"d4e" => DATA <= x"4449";
            when "01" & x"d4f" => DATA <= x"2000";
            when "01" & x"d50" => DATA <= x"003f";
            when "01" & x"d51" => DATA <= x"39e0";
            when "01" & x"d52" => DATA <= x"0a00";
            when "01" & x"d53" => DATA <= x"ff00";
            when "01" & x"d54" => DATA <= x"454f";
            when "01" & x"d55" => DATA <= x"5249";
            when "01" & x"d56" => DATA <= x"2000";
            when "01" & x"d57" => DATA <= x"003f";
            when "01" & x"d58" => DATA <= x"39e0";
            when "01" & x"d59" => DATA <= x"0c00";
            when "01" & x"d5a" => DATA <= x"ff00";
            when "01" & x"d5b" => DATA <= x"434d";
            when "01" & x"d5c" => DATA <= x"5049";
            when "01" & x"d5d" => DATA <= x"2000";
            when "01" & x"d5e" => DATA <= x"003f";
            when "01" & x"d5f" => DATA <= x"39e0";
            when "01" & x"d60" => DATA <= x"0108";
            when "01" & x"d61" => DATA <= x"f138";
            when "01" & x"d62" => DATA <= x"4d4f";
            when "01" & x"d63" => DATA <= x"5645";
            when "01" & x"d64" => DATA <= x"5000";
            when "01" & x"d65" => DATA <= x"003f";
            when "01" & x"d66" => DATA <= x"39e0";
            when "01" & x"d67" => DATA <= x"0100";
            when "01" & x"d68" => DATA <= x"f1c0";
            when "01" & x"d69" => DATA <= x"4254";
            when "01" & x"d6a" => DATA <= x"5354";
            when "01" & x"d6b" => DATA <= x"2000";
            when "01" & x"d6c" => DATA <= x"003f";
            when "01" & x"d6d" => DATA <= x"39e0";
            when "01" & x"d6e" => DATA <= x"0140";
            when "01" & x"d6f" => DATA <= x"f1c0";
            when "01" & x"d70" => DATA <= x"4243";
            when "01" & x"d71" => DATA <= x"4847";
            when "01" & x"d72" => DATA <= x"2000";
            when "01" & x"d73" => DATA <= x"003f";
            when "01" & x"d74" => DATA <= x"39e0";
            when "01" & x"d75" => DATA <= x"0180";
            when "01" & x"d76" => DATA <= x"f1c0";
            when "01" & x"d77" => DATA <= x"4243";
            when "01" & x"d78" => DATA <= x"4c52";
            when "01" & x"d79" => DATA <= x"2000";
            when "01" & x"d7a" => DATA <= x"003f";
            when "01" & x"d7b" => DATA <= x"39e0";
            when "01" & x"d7c" => DATA <= x"01c0";
            when "01" & x"d7d" => DATA <= x"f1c0";
            when "01" & x"d7e" => DATA <= x"4253";
            when "01" & x"d7f" => DATA <= x"4554";
            when "01" & x"d80" => DATA <= x"2000";
            when "01" & x"d81" => DATA <= x"003f";
            when "01" & x"d82" => DATA <= x"39e0";
            when "01" & x"d83" => DATA <= x"0040";
            when "01" & x"d84" => DATA <= x"c1c0";
            when "01" & x"d85" => DATA <= x"4d4f";
            when "01" & x"d86" => DATA <= x"5645";
            when "01" & x"d87" => DATA <= x"4100";
            when "01" & x"d88" => DATA <= x"003f";
            when "01" & x"d89" => DATA <= x"39e0";
            when "01" & x"d8a" => DATA <= x"0000";
            when "01" & x"d8b" => DATA <= x"c000";
            when "01" & x"d8c" => DATA <= x"4d4f";
            when "01" & x"d8d" => DATA <= x"5645";
            when "01" & x"d8e" => DATA <= x"2000";
            when "01" & x"d8f" => DATA <= x"003f";
            when "01" & x"d90" => DATA <= x"39e0";
            when "01" & x"d91" => DATA <= x"4afc";
            when "01" & x"d92" => DATA <= x"ffff";
            when "01" & x"d93" => DATA <= x"494c";
            when "01" & x"d94" => DATA <= x"4c45";
            when "01" & x"d95" => DATA <= x"4700";
            when "01" & x"d96" => DATA <= x"003f";
            when "01" & x"d97" => DATA <= x"39e0";
            when "01" & x"d98" => DATA <= x"4e70";
            when "01" & x"d99" => DATA <= x"ffff";
            when "01" & x"d9a" => DATA <= x"5245";
            when "01" & x"d9b" => DATA <= x"5345";
            when "01" & x"d9c" => DATA <= x"5400";
            when "01" & x"d9d" => DATA <= x"003f";
            when "01" & x"d9e" => DATA <= x"39e0";
            when "01" & x"d9f" => DATA <= x"4e71";
            when "01" & x"da0" => DATA <= x"ffff";
            when "01" & x"da1" => DATA <= x"4e4f";
            when "01" & x"da2" => DATA <= x"5020";
            when "01" & x"da3" => DATA <= x"2000";
            when "01" & x"da4" => DATA <= x"003f";
            when "01" & x"da5" => DATA <= x"39e0";
            when "01" & x"da6" => DATA <= x"4e72";
            when "01" & x"da7" => DATA <= x"ffff";
            when "01" & x"da8" => DATA <= x"5354";
            when "01" & x"da9" => DATA <= x"4f50";
            when "01" & x"daa" => DATA <= x"2000";
            when "01" & x"dab" => DATA <= x"003f";
            when "01" & x"dac" => DATA <= x"39e0";
            when "01" & x"dad" => DATA <= x"4e73";
            when "01" & x"dae" => DATA <= x"ffff";
            when "01" & x"daf" => DATA <= x"5254";
            when "01" & x"db0" => DATA <= x"4520";
            when "01" & x"db1" => DATA <= x"2000";
            when "01" & x"db2" => DATA <= x"003f";
            when "01" & x"db3" => DATA <= x"39e0";
            when "01" & x"db4" => DATA <= x"4e75";
            when "01" & x"db5" => DATA <= x"ffff";
            when "01" & x"db6" => DATA <= x"5254";
            when "01" & x"db7" => DATA <= x"5320";
            when "01" & x"db8" => DATA <= x"2000";
            when "01" & x"db9" => DATA <= x"003f";
            when "01" & x"dba" => DATA <= x"39e0";
            when "01" & x"dbb" => DATA <= x"4e76";
            when "01" & x"dbc" => DATA <= x"ffff";
            when "01" & x"dbd" => DATA <= x"5452";
            when "01" & x"dbe" => DATA <= x"4150";
            when "01" & x"dbf" => DATA <= x"5600";
            when "01" & x"dc0" => DATA <= x"003f";
            when "01" & x"dc1" => DATA <= x"39e0";
            when "01" & x"dc2" => DATA <= x"4e77";
            when "01" & x"dc3" => DATA <= x"ffff";
            when "01" & x"dc4" => DATA <= x"5254";
            when "01" & x"dc5" => DATA <= x"5220";
            when "01" & x"dc6" => DATA <= x"2000";
            when "01" & x"dc7" => DATA <= x"003f";
            when "01" & x"dc8" => DATA <= x"39e0";
            when "01" & x"dc9" => DATA <= x"4840";
            when "01" & x"dca" => DATA <= x"fff8";
            when "01" & x"dcb" => DATA <= x"5357";
            when "01" & x"dcc" => DATA <= x"4150";
            when "01" & x"dcd" => DATA <= x"2000";
            when "01" & x"dce" => DATA <= x"003f";
            when "01" & x"dcf" => DATA <= x"39e0";
            when "01" & x"dd0" => DATA <= x"4e50";
            when "01" & x"dd1" => DATA <= x"fff8";
            when "01" & x"dd2" => DATA <= x"4c49";
            when "01" & x"dd3" => DATA <= x"4e4b";
            when "01" & x"dd4" => DATA <= x"2000";
            when "01" & x"dd5" => DATA <= x"003f";
            when "01" & x"dd6" => DATA <= x"39e0";
            when "01" & x"dd7" => DATA <= x"4e58";
            when "01" & x"dd8" => DATA <= x"fff8";
            when "01" & x"dd9" => DATA <= x"554e";
            when "01" & x"dda" => DATA <= x"4c4b";
            when "01" & x"ddb" => DATA <= x"2000";
            when "01" & x"ddc" => DATA <= x"003f";
            when "01" & x"ddd" => DATA <= x"39e0";
            when "01" & x"dde" => DATA <= x"4e60";
            when "01" & x"ddf" => DATA <= x"fff0";
            when "01" & x"de0" => DATA <= x"4d4f";
            when "01" & x"de1" => DATA <= x"5645";
            when "01" & x"de2" => DATA <= x"2000";
            when "01" & x"de3" => DATA <= x"003f";
            when "01" & x"de4" => DATA <= x"39e0";
            when "01" & x"de5" => DATA <= x"4e40";
            when "01" & x"de6" => DATA <= x"fff0";
            when "01" & x"de7" => DATA <= x"5452";
            when "01" & x"de8" => DATA <= x"4150";
            when "01" & x"de9" => DATA <= x"2000";
            when "01" & x"dea" => DATA <= x"003f";
            when "01" & x"deb" => DATA <= x"39e0";
            when "01" & x"dec" => DATA <= x"4e80";
            when "01" & x"ded" => DATA <= x"ffc0";
            when "01" & x"dee" => DATA <= x"4a53";
            when "01" & x"def" => DATA <= x"5220";
            when "01" & x"df0" => DATA <= x"2000";
            when "01" & x"df1" => DATA <= x"003f";
            when "01" & x"df2" => DATA <= x"39e0";
            when "01" & x"df3" => DATA <= x"4ec0";
            when "01" & x"df4" => DATA <= x"ffc0";
            when "01" & x"df5" => DATA <= x"4a4d";
            when "01" & x"df6" => DATA <= x"5020";
            when "01" & x"df7" => DATA <= x"2000";
            when "01" & x"df8" => DATA <= x"003f";
            when "01" & x"df9" => DATA <= x"39e0";
            when "01" & x"dfa" => DATA <= x"4880";
            when "01" & x"dfb" => DATA <= x"feb8";
            when "01" & x"dfc" => DATA <= x"4558";
            when "01" & x"dfd" => DATA <= x"5420";
            when "01" & x"dfe" => DATA <= x"2000";
            when "01" & x"dff" => DATA <= x"003f";
            when "01" & x"e00" => DATA <= x"39e0";
            when "01" & x"e01" => DATA <= x"40c0";
            when "01" & x"e02" => DATA <= x"ffc0";
            when "01" & x"e03" => DATA <= x"4d4f";
            when "01" & x"e04" => DATA <= x"5645";
            when "01" & x"e05" => DATA <= x"2000";
            when "01" & x"e06" => DATA <= x"003f";
            when "01" & x"e07" => DATA <= x"39e0";
            when "01" & x"e08" => DATA <= x"44c0";
            when "01" & x"e09" => DATA <= x"ffc0";
            when "01" & x"e0a" => DATA <= x"4d4f";
            when "01" & x"e0b" => DATA <= x"5645";
            when "01" & x"e0c" => DATA <= x"2000";
            when "01" & x"e0d" => DATA <= x"003f";
            when "01" & x"e0e" => DATA <= x"39e0";
            when "01" & x"e0f" => DATA <= x"46c0";
            when "01" & x"e10" => DATA <= x"ffc0";
            when "01" & x"e11" => DATA <= x"4d4f";
            when "01" & x"e12" => DATA <= x"5645";
            when "01" & x"e13" => DATA <= x"2000";
            when "01" & x"e14" => DATA <= x"003f";
            when "01" & x"e15" => DATA <= x"39e0";
            when "01" & x"e16" => DATA <= x"4800";
            when "01" & x"e17" => DATA <= x"ffc0";
            when "01" & x"e18" => DATA <= x"4e42";
            when "01" & x"e19" => DATA <= x"4344";
            when "01" & x"e1a" => DATA <= x"2000";
            when "01" & x"e1b" => DATA <= x"003f";
            when "01" & x"e1c" => DATA <= x"39e0";
            when "01" & x"e1d" => DATA <= x"4840";
            when "01" & x"e1e" => DATA <= x"ffc0";
            when "01" & x"e1f" => DATA <= x"5045";
            when "01" & x"e20" => DATA <= x"4120";
            when "01" & x"e21" => DATA <= x"2000";
            when "01" & x"e22" => DATA <= x"003f";
            when "01" & x"e23" => DATA <= x"39e0";
            when "01" & x"e24" => DATA <= x"4ac0";
            when "01" & x"e25" => DATA <= x"ffc0";
            when "01" & x"e26" => DATA <= x"5441";
            when "01" & x"e27" => DATA <= x"5320";
            when "01" & x"e28" => DATA <= x"2000";
            when "01" & x"e29" => DATA <= x"003f";
            when "01" & x"e2a" => DATA <= x"39e0";
            when "01" & x"e2b" => DATA <= x"4000";
            when "01" & x"e2c" => DATA <= x"ff00";
            when "01" & x"e2d" => DATA <= x"4e45";
            when "01" & x"e2e" => DATA <= x"4758";
            when "01" & x"e2f" => DATA <= x"2000";
            when "01" & x"e30" => DATA <= x"003f";
            when "01" & x"e31" => DATA <= x"39e0";
            when "01" & x"e32" => DATA <= x"4200";
            when "01" & x"e33" => DATA <= x"ff00";
            when "01" & x"e34" => DATA <= x"434c";
            when "01" & x"e35" => DATA <= x"5220";
            when "01" & x"e36" => DATA <= x"2000";
            when "01" & x"e37" => DATA <= x"003f";
            when "01" & x"e38" => DATA <= x"39e0";
            when "01" & x"e39" => DATA <= x"4400";
            when "01" & x"e3a" => DATA <= x"ff00";
            when "01" & x"e3b" => DATA <= x"4e45";
            when "01" & x"e3c" => DATA <= x"4720";
            when "01" & x"e3d" => DATA <= x"2000";
            when "01" & x"e3e" => DATA <= x"003f";
            when "01" & x"e3f" => DATA <= x"39e0";
            when "01" & x"e40" => DATA <= x"4600";
            when "01" & x"e41" => DATA <= x"ff00";
            when "01" & x"e42" => DATA <= x"4e4f";
            when "01" & x"e43" => DATA <= x"5420";
            when "01" & x"e44" => DATA <= x"2000";
            when "01" & x"e45" => DATA <= x"003f";
            when "01" & x"e46" => DATA <= x"39e0";
            when "01" & x"e47" => DATA <= x"4a00";
            when "01" & x"e48" => DATA <= x"ff00";
            when "01" & x"e49" => DATA <= x"5453";
            when "01" & x"e4a" => DATA <= x"5420";
            when "01" & x"e4b" => DATA <= x"2000";
            when "01" & x"e4c" => DATA <= x"003f";
            when "01" & x"e4d" => DATA <= x"39e0";
            when "01" & x"e4e" => DATA <= x"4880";
            when "01" & x"e4f" => DATA <= x"fb80";
            when "01" & x"e50" => DATA <= x"4d4f";
            when "01" & x"e51" => DATA <= x"5645";
            when "01" & x"e52" => DATA <= x"4d00";
            when "01" & x"e53" => DATA <= x"003f";
            when "01" & x"e54" => DATA <= x"39e0";
            when "01" & x"e55" => DATA <= x"41c0";
            when "01" & x"e56" => DATA <= x"f1c0";
            when "01" & x"e57" => DATA <= x"4c45";
            when "01" & x"e58" => DATA <= x"4120";
            when "01" & x"e59" => DATA <= x"2000";
            when "01" & x"e5a" => DATA <= x"003f";
            when "01" & x"e5b" => DATA <= x"39e0";
            when "01" & x"e5c" => DATA <= x"4000";
            when "01" & x"e5d" => DATA <= x"f040";
            when "01" & x"e5e" => DATA <= x"4348";
            when "01" & x"e5f" => DATA <= x"4b20";
            when "01" & x"e60" => DATA <= x"2000";
            when "01" & x"e61" => DATA <= x"003f";
            when "01" & x"e62" => DATA <= x"39e0";
            when "01" & x"e63" => DATA <= x"50c8";
            when "01" & x"e64" => DATA <= x"f0f8";
            when "01" & x"e65" => DATA <= x"4442";
            when "01" & x"e66" => DATA <= x"2020";
            when "01" & x"e67" => DATA <= x"2000";
            when "01" & x"e68" => DATA <= x"003f";
            when "01" & x"e69" => DATA <= x"39e0";
            when "01" & x"e6a" => DATA <= x"50c0";
            when "01" & x"e6b" => DATA <= x"f0c0";
            when "01" & x"e6c" => DATA <= x"5320";
            when "01" & x"e6d" => DATA <= x"2020";
            when "01" & x"e6e" => DATA <= x"2000";
            when "01" & x"e6f" => DATA <= x"003f";
            when "01" & x"e70" => DATA <= x"39e0";
            when "01" & x"e71" => DATA <= x"5000";
            when "01" & x"e72" => DATA <= x"f100";
            when "01" & x"e73" => DATA <= x"4144";
            when "01" & x"e74" => DATA <= x"4451";
            when "01" & x"e75" => DATA <= x"2000";
            when "01" & x"e76" => DATA <= x"003f";
            when "01" & x"e77" => DATA <= x"39e0";
            when "01" & x"e78" => DATA <= x"5100";
            when "01" & x"e79" => DATA <= x"f100";
            when "01" & x"e7a" => DATA <= x"5355";
            when "01" & x"e7b" => DATA <= x"4251";
            when "01" & x"e7c" => DATA <= x"2000";
            when "01" & x"e7d" => DATA <= x"003f";
            when "01" & x"e7e" => DATA <= x"39e0";
            when "01" & x"e7f" => DATA <= x"6000";
            when "01" & x"e80" => DATA <= x"ff00";
            when "01" & x"e81" => DATA <= x"4252";
            when "01" & x"e82" => DATA <= x"4120";
            when "01" & x"e83" => DATA <= x"2000";
            when "01" & x"e84" => DATA <= x"003f";
            when "01" & x"e85" => DATA <= x"39e0";
            when "01" & x"e86" => DATA <= x"6100";
            when "01" & x"e87" => DATA <= x"ff00";
            when "01" & x"e88" => DATA <= x"4253";
            when "01" & x"e89" => DATA <= x"5220";
            when "01" & x"e8a" => DATA <= x"2000";
            when "01" & x"e8b" => DATA <= x"003f";
            when "01" & x"e8c" => DATA <= x"39e0";
            when "01" & x"e8d" => DATA <= x"6000";
            when "01" & x"e8e" => DATA <= x"f000";
            when "01" & x"e8f" => DATA <= x"4200";
            when "01" & x"e90" => DATA <= x"0000";
            when "01" & x"e91" => DATA <= x"0000";
            when "01" & x"e92" => DATA <= x"003f";
            when "01" & x"e93" => DATA <= x"39e0";
            when "01" & x"e94" => DATA <= x"7000";
            when "01" & x"e95" => DATA <= x"f100";
            when "01" & x"e96" => DATA <= x"4d4f";
            when "01" & x"e97" => DATA <= x"5645";
            when "01" & x"e98" => DATA <= x"5100";
            when "01" & x"e99" => DATA <= x"003f";
            when "01" & x"e9a" => DATA <= x"39e0";
            when "01" & x"e9b" => DATA <= x"8100";
            when "01" & x"e9c" => DATA <= x"f1f0";
            when "01" & x"e9d" => DATA <= x"5342";
            when "01" & x"e9e" => DATA <= x"4344";
            when "01" & x"e9f" => DATA <= x"2000";
            when "01" & x"ea0" => DATA <= x"003f";
            when "01" & x"ea1" => DATA <= x"39e0";
            when "01" & x"ea2" => DATA <= x"80c0";
            when "01" & x"ea3" => DATA <= x"f1c0";
            when "01" & x"ea4" => DATA <= x"4449";
            when "01" & x"ea5" => DATA <= x"5655";
            when "01" & x"ea6" => DATA <= x"2000";
            when "01" & x"ea7" => DATA <= x"003f";
            when "01" & x"ea8" => DATA <= x"39e0";
            when "01" & x"ea9" => DATA <= x"81c0";
            when "01" & x"eaa" => DATA <= x"f1c0";
            when "01" & x"eab" => DATA <= x"4449";
            when "01" & x"eac" => DATA <= x"5653";
            when "01" & x"ead" => DATA <= x"2000";
            when "01" & x"eae" => DATA <= x"003f";
            when "01" & x"eaf" => DATA <= x"39e0";
            when "01" & x"eb0" => DATA <= x"8000";
            when "01" & x"eb1" => DATA <= x"f000";
            when "01" & x"eb2" => DATA <= x"4f52";
            when "01" & x"eb3" => DATA <= x"2020";
            when "01" & x"eb4" => DATA <= x"2000";
            when "01" & x"eb5" => DATA <= x"003f";
            when "01" & x"eb6" => DATA <= x"39e0";
            when "01" & x"eb7" => DATA <= x"9100";
            when "01" & x"eb8" => DATA <= x"f130";
            when "01" & x"eb9" => DATA <= x"5355";
            when "01" & x"eba" => DATA <= x"4258";
            when "01" & x"ebb" => DATA <= x"2000";
            when "01" & x"ebc" => DATA <= x"003f";
            when "01" & x"ebd" => DATA <= x"39e0";
            when "01" & x"ebe" => DATA <= x"90c0";
            when "01" & x"ebf" => DATA <= x"f0c0";
            when "01" & x"ec0" => DATA <= x"5355";
            when "01" & x"ec1" => DATA <= x"4241";
            when "01" & x"ec2" => DATA <= x"2000";
            when "01" & x"ec3" => DATA <= x"003f";
            when "01" & x"ec4" => DATA <= x"39e0";
            when "01" & x"ec5" => DATA <= x"9000";
            when "01" & x"ec6" => DATA <= x"f000";
            when "01" & x"ec7" => DATA <= x"5355";
            when "01" & x"ec8" => DATA <= x"4220";
            when "01" & x"ec9" => DATA <= x"2000";
            when "01" & x"eca" => DATA <= x"003f";
            when "01" & x"ecb" => DATA <= x"39e0";
            when "01" & x"ecc" => DATA <= x"b108";
            when "01" & x"ecd" => DATA <= x"f138";
            when "01" & x"ece" => DATA <= x"434d";
            when "01" & x"ecf" => DATA <= x"504d";
            when "01" & x"ed0" => DATA <= x"2000";
            when "01" & x"ed1" => DATA <= x"003f";
            when "01" & x"ed2" => DATA <= x"39e0";
            when "01" & x"ed3" => DATA <= x"b0c0";
            when "01" & x"ed4" => DATA <= x"f0c0";
            when "01" & x"ed5" => DATA <= x"434d";
            when "01" & x"ed6" => DATA <= x"5041";
            when "01" & x"ed7" => DATA <= x"2000";
            when "01" & x"ed8" => DATA <= x"003f";
            when "01" & x"ed9" => DATA <= x"39e0";
            when "01" & x"eda" => DATA <= x"b100";
            when "01" & x"edb" => DATA <= x"f100";
            when "01" & x"edc" => DATA <= x"454f";
            when "01" & x"edd" => DATA <= x"5220";
            when "01" & x"ede" => DATA <= x"2000";
            when "01" & x"edf" => DATA <= x"003f";
            when "01" & x"ee0" => DATA <= x"39e0";
            when "01" & x"ee1" => DATA <= x"b000";
            when "01" & x"ee2" => DATA <= x"f000";
            when "01" & x"ee3" => DATA <= x"434d";
            when "01" & x"ee4" => DATA <= x"5020";
            when "01" & x"ee5" => DATA <= x"2000";
            when "01" & x"ee6" => DATA <= x"003f";
            when "01" & x"ee7" => DATA <= x"39e0";
            when "01" & x"ee8" => DATA <= x"c140";
            when "01" & x"ee9" => DATA <= x"f1f8";
            when "01" & x"eea" => DATA <= x"4558";
            when "01" & x"eeb" => DATA <= x"4720";
            when "01" & x"eec" => DATA <= x"2000";
            when "01" & x"eed" => DATA <= x"003f";
            when "01" & x"eee" => DATA <= x"39e0";
            when "01" & x"eef" => DATA <= x"c148";
            when "01" & x"ef0" => DATA <= x"f1f8";
            when "01" & x"ef1" => DATA <= x"4558";
            when "01" & x"ef2" => DATA <= x"4720";
            when "01" & x"ef3" => DATA <= x"2000";
            when "01" & x"ef4" => DATA <= x"003f";
            when "01" & x"ef5" => DATA <= x"39e0";
            when "01" & x"ef6" => DATA <= x"c188";
            when "01" & x"ef7" => DATA <= x"f1f8";
            when "01" & x"ef8" => DATA <= x"4558";
            when "01" & x"ef9" => DATA <= x"4720";
            when "01" & x"efa" => DATA <= x"2000";
            when "01" & x"efb" => DATA <= x"003f";
            when "01" & x"efc" => DATA <= x"39e0";
            when "01" & x"efd" => DATA <= x"c100";
            when "01" & x"efe" => DATA <= x"f1f0";
            when "01" & x"eff" => DATA <= x"4142";
            when "01" & x"f00" => DATA <= x"4344";
            when "01" & x"f01" => DATA <= x"2000";
            when "01" & x"f02" => DATA <= x"003f";
            when "01" & x"f03" => DATA <= x"39e0";
            when "01" & x"f04" => DATA <= x"c1c0";
            when "01" & x"f05" => DATA <= x"f1c0";
            when "01" & x"f06" => DATA <= x"4d55";
            when "01" & x"f07" => DATA <= x"4c53";
            when "01" & x"f08" => DATA <= x"2000";
            when "01" & x"f09" => DATA <= x"003f";
            when "01" & x"f0a" => DATA <= x"39e0";
            when "01" & x"f0b" => DATA <= x"c0c0";
            when "01" & x"f0c" => DATA <= x"f1c0";
            when "01" & x"f0d" => DATA <= x"4d55";
            when "01" & x"f0e" => DATA <= x"4c55";
            when "01" & x"f0f" => DATA <= x"2000";
            when "01" & x"f10" => DATA <= x"003f";
            when "01" & x"f11" => DATA <= x"39e0";
            when "01" & x"f12" => DATA <= x"c000";
            when "01" & x"f13" => DATA <= x"f000";
            when "01" & x"f14" => DATA <= x"414e";
            when "01" & x"f15" => DATA <= x"4420";
            when "01" & x"f16" => DATA <= x"2000";
            when "01" & x"f17" => DATA <= x"003f";
            when "01" & x"f18" => DATA <= x"39e0";
            when "01" & x"f19" => DATA <= x"d100";
            when "01" & x"f1a" => DATA <= x"f130";
            when "01" & x"f1b" => DATA <= x"4144";
            when "01" & x"f1c" => DATA <= x"4458";
            when "01" & x"f1d" => DATA <= x"2000";
            when "01" & x"f1e" => DATA <= x"003f";
            when "01" & x"f1f" => DATA <= x"39e0";
            when "01" & x"f20" => DATA <= x"d0c0";
            when "01" & x"f21" => DATA <= x"f0c0";
            when "01" & x"f22" => DATA <= x"4144";
            when "01" & x"f23" => DATA <= x"4441";
            when "01" & x"f24" => DATA <= x"2000";
            when "01" & x"f25" => DATA <= x"003f";
            when "01" & x"f26" => DATA <= x"39e0";
            when "01" & x"f27" => DATA <= x"d000";
            when "01" & x"f28" => DATA <= x"f000";
            when "01" & x"f29" => DATA <= x"4144";
            when "01" & x"f2a" => DATA <= x"4420";
            when "01" & x"f2b" => DATA <= x"2000";
            when "01" & x"f2c" => DATA <= x"003f";
            when "01" & x"f2d" => DATA <= x"39e0";
            when "01" & x"f2e" => DATA <= x"e0c0";
            when "01" & x"f2f" => DATA <= x"fec0";
            when "01" & x"f30" => DATA <= x"4153";
            when "01" & x"f31" => DATA <= x"2020";
            when "01" & x"f32" => DATA <= x"2000";
            when "01" & x"f33" => DATA <= x"003f";
            when "01" & x"f34" => DATA <= x"39e0";
            when "01" & x"f35" => DATA <= x"e2c0";
            when "01" & x"f36" => DATA <= x"fec0";
            when "01" & x"f37" => DATA <= x"4c53";
            when "01" & x"f38" => DATA <= x"2020";
            when "01" & x"f39" => DATA <= x"2000";
            when "01" & x"f3a" => DATA <= x"003f";
            when "01" & x"f3b" => DATA <= x"39e0";
            when "01" & x"f3c" => DATA <= x"e4c0";
            when "01" & x"f3d" => DATA <= x"fec0";
            when "01" & x"f3e" => DATA <= x"524f";
            when "01" & x"f3f" => DATA <= x"5820";
            when "01" & x"f40" => DATA <= x"2000";
            when "01" & x"f41" => DATA <= x"003f";
            when "01" & x"f42" => DATA <= x"39e0";
            when "01" & x"f43" => DATA <= x"e6c0";
            when "01" & x"f44" => DATA <= x"fec0";
            when "01" & x"f45" => DATA <= x"524f";
            when "01" & x"f46" => DATA <= x"2020";
            when "01" & x"f47" => DATA <= x"2000";
            when "01" & x"f48" => DATA <= x"003f";
            when "01" & x"f49" => DATA <= x"39e0";
            when "01" & x"f4a" => DATA <= x"e000";
            when "01" & x"f4b" => DATA <= x"f018";
            when "01" & x"f4c" => DATA <= x"4153";
            when "01" & x"f4d" => DATA <= x"2020";
            when "01" & x"f4e" => DATA <= x"2000";
            when "01" & x"f4f" => DATA <= x"003f";
            when "01" & x"f50" => DATA <= x"39e0";
            when "01" & x"f51" => DATA <= x"e008";
            when "01" & x"f52" => DATA <= x"f018";
            when "01" & x"f53" => DATA <= x"4c53";
            when "01" & x"f54" => DATA <= x"2020";
            when "01" & x"f55" => DATA <= x"2000";
            when "01" & x"f56" => DATA <= x"003f";
            when "01" & x"f57" => DATA <= x"39e0";
            when "01" & x"f58" => DATA <= x"e010";
            when "01" & x"f59" => DATA <= x"f018";
            when "01" & x"f5a" => DATA <= x"524f";
            when "01" & x"f5b" => DATA <= x"5820";
            when "01" & x"f5c" => DATA <= x"2000";
            when "01" & x"f5d" => DATA <= x"003f";
            when "01" & x"f5e" => DATA <= x"39e0";
            when "01" & x"f5f" => DATA <= x"e018";
            when "01" & x"f60" => DATA <= x"f018";
            when "01" & x"f61" => DATA <= x"524f";
            when "01" & x"f62" => DATA <= x"2020";
            when "01" & x"f63" => DATA <= x"2000";
            when "01" & x"f64" => DATA <= x"003f";
            when "01" & x"f65" => DATA <= x"39e0";
            when "01" & x"f66" => DATA <= x"0000";
            when "01" & x"f67" => DATA <= x"0000";
            when "01" & x"f68" => DATA <= x"3f3f";
            when "01" & x"f69" => DATA <= x"3f3f";
            when "01" & x"f6a" => DATA <= x"3f00";
            when "01" & x"f6b" => DATA <= x"003f";
            when "01" & x"f6c" => DATA <= x"39e0";
            when "01" & x"f6d" => DATA <= x"2532";
            when "01" & x"f6e" => DATA <= x"343a";
            when "01" & x"f6f" => DATA <= x"256d";
            when "01" & x"f70" => DATA <= x"693a";
            when "01" & x"f71" => DATA <= x"2573";
            when "01" & x"f72" => DATA <= x"6520";
            when "01" & x"f73" => DATA <= x"2564";
            when "01" & x"f74" => DATA <= x"792d";
            when "01" & x"f75" => DATA <= x"256d";
            when "01" & x"f76" => DATA <= x"332d";
            when "01" & x"f77" => DATA <= x"2563";
            when "01" & x"f78" => DATA <= x"6525";
            when "01" & x"f79" => DATA <= x"7972";
            when "01" & x"f7a" => DATA <= x"0006";
            when "01" & x"f7b" => DATA <= x"7c00";
            when "01" & x"f7c" => DATA <= x"5206";
            when "01" & x"f7d" => DATA <= x"bcbc";
            when "01" & x"f7e" => DATA <= x"0010";
            when "01" & x"f7f" => DATA <= x"0000";
            when "01" & x"f80" => DATA <= x"66f6";
            when "01" & x"f81" => DATA <= x"103c";
            when "01" & x"f82" => DATA <= x"002a";
            when "01" & x"f83" => DATA <= x"6100";
            when "01" & x"f84" => DATA <= x"cade";
            when "01" & x"f85" => DATA <= x"60e9";
            when "01" & x"f86" => DATA <= x"002a";
            when "01" & x"f87" => DATA <= x"6100";
            when "01" & x"f88" => DATA <= x"cae0";
            when "01" & x"f89" => DATA <= x"60e9";
            when "01" & x"f8a" => DATA <= x"cade";
            when "01" & x"f8b" => DATA <= x"60e9";
            when "01" & x"f8c" => DATA <= x"ffff";
            when "01" & x"f8d" => DATA <= x"ffff";
            when "01" & x"f8e" => DATA <= x"ffff";
            when "01" & x"f8f" => DATA <= x"ffff";
            when "01" & x"f90" => DATA <= x"ffff";
            when "01" & x"f91" => DATA <= x"ffff";
            when "01" & x"f92" => DATA <= x"ffff";
            when "01" & x"f93" => DATA <= x"ffff";
            when "01" & x"f94" => DATA <= x"ffff";
            when "01" & x"f95" => DATA <= x"ffff";
            when "01" & x"f96" => DATA <= x"ffff";
            when "01" & x"f97" => DATA <= x"ffff";
            when "01" & x"f98" => DATA <= x"ffff";
            when "01" & x"f99" => DATA <= x"ffff";
            when "01" & x"f9a" => DATA <= x"ffff";
            when "01" & x"f9b" => DATA <= x"ffff";
            when "01" & x"f9c" => DATA <= x"ffff";
            when "01" & x"f9d" => DATA <= x"ffff";
            when "01" & x"f9e" => DATA <= x"ffff";
            when "01" & x"f9f" => DATA <= x"ffff";
            when "01" & x"fa0" => DATA <= x"ffff";
            when "01" & x"fa1" => DATA <= x"ffff";
            when "01" & x"fa2" => DATA <= x"ffff";
            when "01" & x"fa3" => DATA <= x"ffff";
            when "01" & x"fa4" => DATA <= x"ffff";
            when "01" & x"fa5" => DATA <= x"ffff";
            when "01" & x"fa6" => DATA <= x"ffff";
            when "01" & x"fa7" => DATA <= x"ffff";
            when "01" & x"fa8" => DATA <= x"ffff";
            when "01" & x"fa9" => DATA <= x"ffff";
            when "01" & x"faa" => DATA <= x"ffff";
            when "01" & x"fab" => DATA <= x"ffff";
            when "01" & x"fac" => DATA <= x"ffff";
            when "01" & x"fad" => DATA <= x"ffff";
            when "01" & x"fae" => DATA <= x"ffff";
            when "01" & x"faf" => DATA <= x"ffff";
            when "01" & x"fb0" => DATA <= x"ffff";
            when "01" & x"fb1" => DATA <= x"ffff";
            when "01" & x"fb2" => DATA <= x"ffff";
            when "01" & x"fb3" => DATA <= x"ffff";
            when "01" & x"fb4" => DATA <= x"ffff";
            when "01" & x"fb5" => DATA <= x"ffff";
            when "01" & x"fb6" => DATA <= x"ffff";
            when "01" & x"fb7" => DATA <= x"ffff";
            when "01" & x"fb8" => DATA <= x"ffff";
            when "01" & x"fb9" => DATA <= x"ffff";
            when "01" & x"fba" => DATA <= x"ffff";
            when "01" & x"fbb" => DATA <= x"ffff";
            when "01" & x"fbc" => DATA <= x"ffff";
            when "01" & x"fbd" => DATA <= x"ffff";
            when "01" & x"fbe" => DATA <= x"ffff";
            when "01" & x"fbf" => DATA <= x"ffff";
            when "01" & x"fc0" => DATA <= x"ffff";
            when "01" & x"fc1" => DATA <= x"ffff";
            when "01" & x"fc2" => DATA <= x"ffff";
            when "01" & x"fc3" => DATA <= x"ffff";
            when "01" & x"fc4" => DATA <= x"ffff";
            when "01" & x"fc5" => DATA <= x"ffff";
            when "01" & x"fc6" => DATA <= x"ffff";
            when "01" & x"fc7" => DATA <= x"ffff";
            when "01" & x"fc8" => DATA <= x"ffff";
            when "01" & x"fc9" => DATA <= x"ffff";
            when "01" & x"fca" => DATA <= x"ffff";
            when "01" & x"fcb" => DATA <= x"ffff";
            when "01" & x"fcc" => DATA <= x"ffff";
            when "01" & x"fcd" => DATA <= x"ffff";
            when "01" & x"fce" => DATA <= x"ffff";
            when "01" & x"fcf" => DATA <= x"ffff";
            when "01" & x"fd0" => DATA <= x"ffff";
            when "01" & x"fd1" => DATA <= x"ffff";
            when "01" & x"fd2" => DATA <= x"ffff";
            when "01" & x"fd3" => DATA <= x"ffff";
            when "01" & x"fd4" => DATA <= x"ffff";
            when "01" & x"fd5" => DATA <= x"ffff";
            when "01" & x"fd6" => DATA <= x"ffff";
            when "01" & x"fd7" => DATA <= x"ffff";
            when "01" & x"fd8" => DATA <= x"ffff";
            when "01" & x"fd9" => DATA <= x"ffff";
            when "01" & x"fda" => DATA <= x"ffff";
            when "01" & x"fdb" => DATA <= x"ffff";
            when "01" & x"fdc" => DATA <= x"ffff";
            when "01" & x"fdd" => DATA <= x"ffff";
            when "01" & x"fde" => DATA <= x"ffff";
            when "01" & x"fdf" => DATA <= x"ffff";
            when "01" & x"fe0" => DATA <= x"ffff";
            when "01" & x"fe1" => DATA <= x"ffff";
            when "01" & x"fe2" => DATA <= x"ffff";
            when "01" & x"fe3" => DATA <= x"ffff";
            when "01" & x"fe4" => DATA <= x"ffff";
            when "01" & x"fe5" => DATA <= x"ffff";
            when "01" & x"fe6" => DATA <= x"ffff";
            when "01" & x"fe7" => DATA <= x"ffff";
            when "01" & x"fe8" => DATA <= x"ffff";
            when "01" & x"fe9" => DATA <= x"ffff";
            when "01" & x"fea" => DATA <= x"ffff";
            when "01" & x"feb" => DATA <= x"ffff";
            when "01" & x"fec" => DATA <= x"ffff";
            when "01" & x"fed" => DATA <= x"ffff";
            when "01" & x"fee" => DATA <= x"ffff";
            when "01" & x"fef" => DATA <= x"ffff";
            when "01" & x"ff0" => DATA <= x"ffff";
            when "01" & x"ff1" => DATA <= x"ffff";
            when "01" & x"ff2" => DATA <= x"ffff";
            when "01" & x"ff3" => DATA <= x"ffff";
            when "01" & x"ff4" => DATA <= x"ffff";
            when "01" & x"ff5" => DATA <= x"ffff";
            when "01" & x"ff6" => DATA <= x"ffff";
            when "01" & x"ff7" => DATA <= x"ffff";
            when "01" & x"ff8" => DATA <= x"ffff";
            when "01" & x"ff9" => DATA <= x"ffff";
            when "01" & x"ffa" => DATA <= x"ffff";
            when "01" & x"ffb" => DATA <= x"ffff";
            when "01" & x"ffc" => DATA <= x"ffff";
            when "01" & x"ffd" => DATA <= x"ffff";
            when "01" & x"ffe" => DATA <= x"ffff";
            when "01" & x"fff" => DATA <= x"ffff";
            when "10" & x"000" => DATA <= x"ffff";
            when "10" & x"001" => DATA <= x"ffff";
            when "10" & x"002" => DATA <= x"ffff";
            when "10" & x"003" => DATA <= x"ffff";
            when "10" & x"004" => DATA <= x"ffff";
            when "10" & x"005" => DATA <= x"ffff";
            when "10" & x"006" => DATA <= x"ffff";
            when "10" & x"007" => DATA <= x"ffff";
            when "10" & x"008" => DATA <= x"ffff";
            when "10" & x"009" => DATA <= x"ffff";
            when "10" & x"00a" => DATA <= x"ffff";
            when "10" & x"00b" => DATA <= x"ffff";
            when "10" & x"00c" => DATA <= x"ffff";
            when "10" & x"00d" => DATA <= x"ffff";
            when "10" & x"00e" => DATA <= x"ffff";
            when "10" & x"00f" => DATA <= x"ffff";
            when "10" & x"010" => DATA <= x"ffff";
            when "10" & x"011" => DATA <= x"ffff";
            when "10" & x"012" => DATA <= x"ffff";
            when "10" & x"013" => DATA <= x"ffff";
            when "10" & x"014" => DATA <= x"ffff";
            when "10" & x"015" => DATA <= x"ffff";
            when "10" & x"016" => DATA <= x"ffff";
            when "10" & x"017" => DATA <= x"ffff";
            when "10" & x"018" => DATA <= x"ffff";
            when "10" & x"019" => DATA <= x"ffff";
            when "10" & x"01a" => DATA <= x"ffff";
            when "10" & x"01b" => DATA <= x"ffff";
            when "10" & x"01c" => DATA <= x"ffff";
            when "10" & x"01d" => DATA <= x"ffff";
            when "10" & x"01e" => DATA <= x"ffff";
            when "10" & x"01f" => DATA <= x"ffff";
            when "10" & x"020" => DATA <= x"ffff";
            when "10" & x"021" => DATA <= x"ffff";
            when "10" & x"022" => DATA <= x"ffff";
            when "10" & x"023" => DATA <= x"ffff";
            when "10" & x"024" => DATA <= x"ffff";
            when "10" & x"025" => DATA <= x"ffff";
            when "10" & x"026" => DATA <= x"ffff";
            when "10" & x"027" => DATA <= x"ffff";
            when "10" & x"028" => DATA <= x"ffff";
            when "10" & x"029" => DATA <= x"ffff";
            when "10" & x"02a" => DATA <= x"ffff";
            when "10" & x"02b" => DATA <= x"ffff";
            when "10" & x"02c" => DATA <= x"ffff";
            when "10" & x"02d" => DATA <= x"ffff";
            when "10" & x"02e" => DATA <= x"ffff";
            when "10" & x"02f" => DATA <= x"ffff";
            when "10" & x"030" => DATA <= x"ffff";
            when "10" & x"031" => DATA <= x"ffff";
            when "10" & x"032" => DATA <= x"ffff";
            when "10" & x"033" => DATA <= x"ffff";
            when "10" & x"034" => DATA <= x"ffff";
            when "10" & x"035" => DATA <= x"ffff";
            when "10" & x"036" => DATA <= x"ffff";
            when "10" & x"037" => DATA <= x"ffff";
            when "10" & x"038" => DATA <= x"ffff";
            when "10" & x"039" => DATA <= x"ffff";
            when "10" & x"03a" => DATA <= x"ffff";
            when "10" & x"03b" => DATA <= x"ffff";
            when "10" & x"03c" => DATA <= x"ffff";
            when "10" & x"03d" => DATA <= x"ffff";
            when "10" & x"03e" => DATA <= x"ffff";
            when "10" & x"03f" => DATA <= x"ffff";
            when "10" & x"040" => DATA <= x"ffff";
            when "10" & x"041" => DATA <= x"ffff";
            when "10" & x"042" => DATA <= x"ffff";
            when "10" & x"043" => DATA <= x"ffff";
            when "10" & x"044" => DATA <= x"ffff";
            when "10" & x"045" => DATA <= x"ffff";
            when "10" & x"046" => DATA <= x"ffff";
            when "10" & x"047" => DATA <= x"ffff";
            when "10" & x"048" => DATA <= x"ffff";
            when "10" & x"049" => DATA <= x"ffff";
            when "10" & x"04a" => DATA <= x"ffff";
            when "10" & x"04b" => DATA <= x"ffff";
            when "10" & x"04c" => DATA <= x"ffff";
            when "10" & x"04d" => DATA <= x"ffff";
            when "10" & x"04e" => DATA <= x"ffff";
            when "10" & x"04f" => DATA <= x"ffff";
            when "10" & x"050" => DATA <= x"ffff";
            when "10" & x"051" => DATA <= x"ffff";
            when "10" & x"052" => DATA <= x"ffff";
            when "10" & x"053" => DATA <= x"ffff";
            when "10" & x"054" => DATA <= x"ffff";
            when "10" & x"055" => DATA <= x"ffff";
            when "10" & x"056" => DATA <= x"ffff";
            when "10" & x"057" => DATA <= x"ffff";
            when "10" & x"058" => DATA <= x"ffff";
            when "10" & x"059" => DATA <= x"ffff";
            when "10" & x"05a" => DATA <= x"ffff";
            when "10" & x"05b" => DATA <= x"ffff";
            when "10" & x"05c" => DATA <= x"ffff";
            when "10" & x"05d" => DATA <= x"ffff";
            when "10" & x"05e" => DATA <= x"ffff";
            when "10" & x"05f" => DATA <= x"ffff";
            when "10" & x"060" => DATA <= x"ffff";
            when "10" & x"061" => DATA <= x"ffff";
            when "10" & x"062" => DATA <= x"ffff";
            when "10" & x"063" => DATA <= x"ffff";
            when "10" & x"064" => DATA <= x"ffff";
            when "10" & x"065" => DATA <= x"ffff";
            when "10" & x"066" => DATA <= x"ffff";
            when "10" & x"067" => DATA <= x"ffff";
            when "10" & x"068" => DATA <= x"ffff";
            when "10" & x"069" => DATA <= x"ffff";
            when "10" & x"06a" => DATA <= x"ffff";
            when "10" & x"06b" => DATA <= x"ffff";
            when "10" & x"06c" => DATA <= x"ffff";
            when "10" & x"06d" => DATA <= x"ffff";
            when "10" & x"06e" => DATA <= x"ffff";
            when "10" & x"06f" => DATA <= x"ffff";
            when "10" & x"070" => DATA <= x"ffff";
            when "10" & x"071" => DATA <= x"ffff";
            when "10" & x"072" => DATA <= x"ffff";
            when "10" & x"073" => DATA <= x"ffff";
            when "10" & x"074" => DATA <= x"ffff";
            when "10" & x"075" => DATA <= x"ffff";
            when "10" & x"076" => DATA <= x"ffff";
            when "10" & x"077" => DATA <= x"ffff";
            when "10" & x"078" => DATA <= x"ffff";
            when "10" & x"079" => DATA <= x"ffff";
            when "10" & x"07a" => DATA <= x"ffff";
            when "10" & x"07b" => DATA <= x"ffff";
            when "10" & x"07c" => DATA <= x"ffff";
            when "10" & x"07d" => DATA <= x"ffff";
            when "10" & x"07e" => DATA <= x"ffff";
            when "10" & x"07f" => DATA <= x"ffff";
            when "10" & x"080" => DATA <= x"ffff";
            when "10" & x"081" => DATA <= x"ffff";
            when "10" & x"082" => DATA <= x"ffff";
            when "10" & x"083" => DATA <= x"ffff";
            when "10" & x"084" => DATA <= x"ffff";
            when "10" & x"085" => DATA <= x"ffff";
            when "10" & x"086" => DATA <= x"ffff";
            when "10" & x"087" => DATA <= x"ffff";
            when "10" & x"088" => DATA <= x"ffff";
            when "10" & x"089" => DATA <= x"ffff";
            when "10" & x"08a" => DATA <= x"ffff";
            when "10" & x"08b" => DATA <= x"ffff";
            when "10" & x"08c" => DATA <= x"ffff";
            when "10" & x"08d" => DATA <= x"ffff";
            when "10" & x"08e" => DATA <= x"ffff";
            when "10" & x"08f" => DATA <= x"ffff";
            when "10" & x"090" => DATA <= x"ffff";
            when "10" & x"091" => DATA <= x"ffff";
            when "10" & x"092" => DATA <= x"ffff";
            when "10" & x"093" => DATA <= x"ffff";
            when "10" & x"094" => DATA <= x"ffff";
            when "10" & x"095" => DATA <= x"ffff";
            when "10" & x"096" => DATA <= x"ffff";
            when "10" & x"097" => DATA <= x"ffff";
            when "10" & x"098" => DATA <= x"ffff";
            when "10" & x"099" => DATA <= x"ffff";
            when "10" & x"09a" => DATA <= x"ffff";
            when "10" & x"09b" => DATA <= x"ffff";
            when "10" & x"09c" => DATA <= x"ffff";
            when "10" & x"09d" => DATA <= x"ffff";
            when "10" & x"09e" => DATA <= x"ffff";
            when "10" & x"09f" => DATA <= x"ffff";
            when "10" & x"0a0" => DATA <= x"ffff";
            when "10" & x"0a1" => DATA <= x"ffff";
            when "10" & x"0a2" => DATA <= x"ffff";
            when "10" & x"0a3" => DATA <= x"ffff";
            when "10" & x"0a4" => DATA <= x"ffff";
            when "10" & x"0a5" => DATA <= x"ffff";
            when "10" & x"0a6" => DATA <= x"ffff";
            when "10" & x"0a7" => DATA <= x"ffff";
            when "10" & x"0a8" => DATA <= x"ffff";
            when "10" & x"0a9" => DATA <= x"ffff";
            when "10" & x"0aa" => DATA <= x"ffff";
            when "10" & x"0ab" => DATA <= x"ffff";
            when "10" & x"0ac" => DATA <= x"ffff";
            when "10" & x"0ad" => DATA <= x"ffff";
            when "10" & x"0ae" => DATA <= x"ffff";
            when "10" & x"0af" => DATA <= x"ffff";
            when "10" & x"0b0" => DATA <= x"ffff";
            when "10" & x"0b1" => DATA <= x"ffff";
            when "10" & x"0b2" => DATA <= x"ffff";
            when "10" & x"0b3" => DATA <= x"ffff";
            when "10" & x"0b4" => DATA <= x"ffff";
            when "10" & x"0b5" => DATA <= x"ffff";
            when "10" & x"0b6" => DATA <= x"ffff";
            when "10" & x"0b7" => DATA <= x"ffff";
            when "10" & x"0b8" => DATA <= x"ffff";
            when "10" & x"0b9" => DATA <= x"ffff";
            when "10" & x"0ba" => DATA <= x"ffff";
            when "10" & x"0bb" => DATA <= x"ffff";
            when "10" & x"0bc" => DATA <= x"ffff";
            when "10" & x"0bd" => DATA <= x"ffff";
            when "10" & x"0be" => DATA <= x"ffff";
            when "10" & x"0bf" => DATA <= x"ffff";
            when "10" & x"0c0" => DATA <= x"ffff";
            when "10" & x"0c1" => DATA <= x"ffff";
            when "10" & x"0c2" => DATA <= x"ffff";
            when "10" & x"0c3" => DATA <= x"ffff";
            when "10" & x"0c4" => DATA <= x"ffff";
            when "10" & x"0c5" => DATA <= x"ffff";
            when "10" & x"0c6" => DATA <= x"ffff";
            when "10" & x"0c7" => DATA <= x"ffff";
            when "10" & x"0c8" => DATA <= x"ffff";
            when "10" & x"0c9" => DATA <= x"ffff";
            when "10" & x"0ca" => DATA <= x"ffff";
            when "10" & x"0cb" => DATA <= x"ffff";
            when "10" & x"0cc" => DATA <= x"ffff";
            when "10" & x"0cd" => DATA <= x"ffff";
            when "10" & x"0ce" => DATA <= x"ffff";
            when "10" & x"0cf" => DATA <= x"ffff";
            when "10" & x"0d0" => DATA <= x"ffff";
            when "10" & x"0d1" => DATA <= x"ffff";
            when "10" & x"0d2" => DATA <= x"ffff";
            when "10" & x"0d3" => DATA <= x"ffff";
            when "10" & x"0d4" => DATA <= x"ffff";
            when "10" & x"0d5" => DATA <= x"ffff";
            when "10" & x"0d6" => DATA <= x"ffff";
            when "10" & x"0d7" => DATA <= x"ffff";
            when "10" & x"0d8" => DATA <= x"ffff";
            when "10" & x"0d9" => DATA <= x"ffff";
            when "10" & x"0da" => DATA <= x"ffff";
            when "10" & x"0db" => DATA <= x"ffff";
            when "10" & x"0dc" => DATA <= x"ffff";
            when "10" & x"0dd" => DATA <= x"ffff";
            when "10" & x"0de" => DATA <= x"ffff";
            when "10" & x"0df" => DATA <= x"ffff";
            when "10" & x"0e0" => DATA <= x"ffff";
            when "10" & x"0e1" => DATA <= x"ffff";
            when "10" & x"0e2" => DATA <= x"ffff";
            when "10" & x"0e3" => DATA <= x"ffff";
            when "10" & x"0e4" => DATA <= x"ffff";
            when "10" & x"0e5" => DATA <= x"ffff";
            when "10" & x"0e6" => DATA <= x"ffff";
            when "10" & x"0e7" => DATA <= x"ffff";
            when "10" & x"0e8" => DATA <= x"ffff";
            when "10" & x"0e9" => DATA <= x"ffff";
            when "10" & x"0ea" => DATA <= x"ffff";
            when "10" & x"0eb" => DATA <= x"ffff";
            when "10" & x"0ec" => DATA <= x"ffff";
            when "10" & x"0ed" => DATA <= x"ffff";
            when "10" & x"0ee" => DATA <= x"ffff";
            when "10" & x"0ef" => DATA <= x"ffff";
            when "10" & x"0f0" => DATA <= x"ffff";
            when "10" & x"0f1" => DATA <= x"ffff";
            when "10" & x"0f2" => DATA <= x"ffff";
            when "10" & x"0f3" => DATA <= x"ffff";
            when "10" & x"0f4" => DATA <= x"ffff";
            when "10" & x"0f5" => DATA <= x"ffff";
            when "10" & x"0f6" => DATA <= x"ffff";
            when "10" & x"0f7" => DATA <= x"ffff";
            when "10" & x"0f8" => DATA <= x"ffff";
            when "10" & x"0f9" => DATA <= x"ffff";
            when "10" & x"0fa" => DATA <= x"ffff";
            when "10" & x"0fb" => DATA <= x"ffff";
            when "10" & x"0fc" => DATA <= x"ffff";
            when "10" & x"0fd" => DATA <= x"ffff";
            when "10" & x"0fe" => DATA <= x"ffff";
            when "10" & x"0ff" => DATA <= x"ffff";
            when "10" & x"100" => DATA <= x"ffff";
            when "10" & x"101" => DATA <= x"ffff";
            when "10" & x"102" => DATA <= x"ffff";
            when "10" & x"103" => DATA <= x"ffff";
            when "10" & x"104" => DATA <= x"ffff";
            when "10" & x"105" => DATA <= x"ffff";
            when "10" & x"106" => DATA <= x"ffff";
            when "10" & x"107" => DATA <= x"ffff";
            when "10" & x"108" => DATA <= x"ffff";
            when "10" & x"109" => DATA <= x"ffff";
            when "10" & x"10a" => DATA <= x"ffff";
            when "10" & x"10b" => DATA <= x"ffff";
            when "10" & x"10c" => DATA <= x"ffff";
            when "10" & x"10d" => DATA <= x"ffff";
            when "10" & x"10e" => DATA <= x"ffff";
            when "10" & x"10f" => DATA <= x"ffff";
            when "10" & x"110" => DATA <= x"ffff";
            when "10" & x"111" => DATA <= x"ffff";
            when "10" & x"112" => DATA <= x"ffff";
            when "10" & x"113" => DATA <= x"ffff";
            when "10" & x"114" => DATA <= x"ffff";
            when "10" & x"115" => DATA <= x"ffff";
            when "10" & x"116" => DATA <= x"ffff";
            when "10" & x"117" => DATA <= x"ffff";
            when "10" & x"118" => DATA <= x"ffff";
            when "10" & x"119" => DATA <= x"ffff";
            when "10" & x"11a" => DATA <= x"ffff";
            when "10" & x"11b" => DATA <= x"ffff";
            when "10" & x"11c" => DATA <= x"ffff";
            when "10" & x"11d" => DATA <= x"ffff";
            when "10" & x"11e" => DATA <= x"ffff";
            when "10" & x"11f" => DATA <= x"ffff";
            when "10" & x"120" => DATA <= x"ffff";
            when "10" & x"121" => DATA <= x"ffff";
            when "10" & x"122" => DATA <= x"ffff";
            when "10" & x"123" => DATA <= x"ffff";
            when "10" & x"124" => DATA <= x"ffff";
            when "10" & x"125" => DATA <= x"ffff";
            when "10" & x"126" => DATA <= x"ffff";
            when "10" & x"127" => DATA <= x"ffff";
            when "10" & x"128" => DATA <= x"ffff";
            when "10" & x"129" => DATA <= x"ffff";
            when "10" & x"12a" => DATA <= x"ffff";
            when "10" & x"12b" => DATA <= x"ffff";
            when "10" & x"12c" => DATA <= x"ffff";
            when "10" & x"12d" => DATA <= x"ffff";
            when "10" & x"12e" => DATA <= x"ffff";
            when "10" & x"12f" => DATA <= x"ffff";
            when "10" & x"130" => DATA <= x"ffff";
            when "10" & x"131" => DATA <= x"ffff";
            when "10" & x"132" => DATA <= x"ffff";
            when "10" & x"133" => DATA <= x"ffff";
            when "10" & x"134" => DATA <= x"ffff";
            when "10" & x"135" => DATA <= x"ffff";
            when "10" & x"136" => DATA <= x"ffff";
            when "10" & x"137" => DATA <= x"ffff";
            when "10" & x"138" => DATA <= x"ffff";
            when "10" & x"139" => DATA <= x"ffff";
            when "10" & x"13a" => DATA <= x"ffff";
            when "10" & x"13b" => DATA <= x"ffff";
            when "10" & x"13c" => DATA <= x"ffff";
            when "10" & x"13d" => DATA <= x"ffff";
            when "10" & x"13e" => DATA <= x"ffff";
            when "10" & x"13f" => DATA <= x"ffff";
            when "10" & x"140" => DATA <= x"ffff";
            when "10" & x"141" => DATA <= x"ffff";
            when "10" & x"142" => DATA <= x"ffff";
            when "10" & x"143" => DATA <= x"ffff";
            when "10" & x"144" => DATA <= x"ffff";
            when "10" & x"145" => DATA <= x"ffff";
            when "10" & x"146" => DATA <= x"ffff";
            when "10" & x"147" => DATA <= x"ffff";
            when "10" & x"148" => DATA <= x"ffff";
            when "10" & x"149" => DATA <= x"ffff";
            when "10" & x"14a" => DATA <= x"ffff";
            when "10" & x"14b" => DATA <= x"ffff";
            when "10" & x"14c" => DATA <= x"ffff";
            when "10" & x"14d" => DATA <= x"ffff";
            when "10" & x"14e" => DATA <= x"ffff";
            when "10" & x"14f" => DATA <= x"ffff";
            when "10" & x"150" => DATA <= x"ffff";
            when "10" & x"151" => DATA <= x"ffff";
            when "10" & x"152" => DATA <= x"ffff";
            when "10" & x"153" => DATA <= x"ffff";
            when "10" & x"154" => DATA <= x"ffff";
            when "10" & x"155" => DATA <= x"ffff";
            when "10" & x"156" => DATA <= x"ffff";
            when "10" & x"157" => DATA <= x"ffff";
            when "10" & x"158" => DATA <= x"ffff";
            when "10" & x"159" => DATA <= x"ffff";
            when "10" & x"15a" => DATA <= x"ffff";
            when "10" & x"15b" => DATA <= x"ffff";
            when "10" & x"15c" => DATA <= x"ffff";
            when "10" & x"15d" => DATA <= x"ffff";
            when "10" & x"15e" => DATA <= x"ffff";
            when "10" & x"15f" => DATA <= x"ffff";
            when "10" & x"160" => DATA <= x"ffff";
            when "10" & x"161" => DATA <= x"ffff";
            when "10" & x"162" => DATA <= x"ffff";
            when "10" & x"163" => DATA <= x"ffff";
            when "10" & x"164" => DATA <= x"ffff";
            when "10" & x"165" => DATA <= x"ffff";
            when "10" & x"166" => DATA <= x"ffff";
            when "10" & x"167" => DATA <= x"ffff";
            when "10" & x"168" => DATA <= x"ffff";
            when "10" & x"169" => DATA <= x"ffff";
            when "10" & x"16a" => DATA <= x"ffff";
            when "10" & x"16b" => DATA <= x"ffff";
            when "10" & x"16c" => DATA <= x"ffff";
            when "10" & x"16d" => DATA <= x"ffff";
            when "10" & x"16e" => DATA <= x"ffff";
            when "10" & x"16f" => DATA <= x"ffff";
            when "10" & x"170" => DATA <= x"ffff";
            when "10" & x"171" => DATA <= x"ffff";
            when "10" & x"172" => DATA <= x"ffff";
            when "10" & x"173" => DATA <= x"ffff";
            when "10" & x"174" => DATA <= x"ffff";
            when "10" & x"175" => DATA <= x"ffff";
            when "10" & x"176" => DATA <= x"ffff";
            when "10" & x"177" => DATA <= x"ffff";
            when "10" & x"178" => DATA <= x"ffff";
            when "10" & x"179" => DATA <= x"ffff";
            when "10" & x"17a" => DATA <= x"ffff";
            when "10" & x"17b" => DATA <= x"ffff";
            when "10" & x"17c" => DATA <= x"ffff";
            when "10" & x"17d" => DATA <= x"ffff";
            when "10" & x"17e" => DATA <= x"ffff";
            when "10" & x"17f" => DATA <= x"ffff";
            when "10" & x"180" => DATA <= x"ffff";
            when "10" & x"181" => DATA <= x"ffff";
            when "10" & x"182" => DATA <= x"ffff";
            when "10" & x"183" => DATA <= x"ffff";
            when "10" & x"184" => DATA <= x"ffff";
            when "10" & x"185" => DATA <= x"ffff";
            when "10" & x"186" => DATA <= x"ffff";
            when "10" & x"187" => DATA <= x"ffff";
            when "10" & x"188" => DATA <= x"ffff";
            when "10" & x"189" => DATA <= x"ffff";
            when "10" & x"18a" => DATA <= x"ffff";
            when "10" & x"18b" => DATA <= x"ffff";
            when "10" & x"18c" => DATA <= x"ffff";
            when "10" & x"18d" => DATA <= x"ffff";
            when "10" & x"18e" => DATA <= x"ffff";
            when "10" & x"18f" => DATA <= x"ffff";
            when "10" & x"190" => DATA <= x"ffff";
            when "10" & x"191" => DATA <= x"ffff";
            when "10" & x"192" => DATA <= x"ffff";
            when "10" & x"193" => DATA <= x"ffff";
            when "10" & x"194" => DATA <= x"ffff";
            when "10" & x"195" => DATA <= x"ffff";
            when "10" & x"196" => DATA <= x"ffff";
            when "10" & x"197" => DATA <= x"ffff";
            when "10" & x"198" => DATA <= x"ffff";
            when "10" & x"199" => DATA <= x"ffff";
            when "10" & x"19a" => DATA <= x"ffff";
            when "10" & x"19b" => DATA <= x"ffff";
            when "10" & x"19c" => DATA <= x"ffff";
            when "10" & x"19d" => DATA <= x"ffff";
            when "10" & x"19e" => DATA <= x"ffff";
            when "10" & x"19f" => DATA <= x"ffff";
            when "10" & x"1a0" => DATA <= x"ffff";
            when "10" & x"1a1" => DATA <= x"ffff";
            when "10" & x"1a2" => DATA <= x"ffff";
            when "10" & x"1a3" => DATA <= x"ffff";
            when "10" & x"1a4" => DATA <= x"ffff";
            when "10" & x"1a5" => DATA <= x"ffff";
            when "10" & x"1a6" => DATA <= x"ffff";
            when "10" & x"1a7" => DATA <= x"ffff";
            when "10" & x"1a8" => DATA <= x"ffff";
            when "10" & x"1a9" => DATA <= x"ffff";
            when "10" & x"1aa" => DATA <= x"ffff";
            when "10" & x"1ab" => DATA <= x"ffff";
            when "10" & x"1ac" => DATA <= x"ffff";
            when "10" & x"1ad" => DATA <= x"ffff";
            when "10" & x"1ae" => DATA <= x"ffff";
            when "10" & x"1af" => DATA <= x"ffff";
            when "10" & x"1b0" => DATA <= x"ffff";
            when "10" & x"1b1" => DATA <= x"ffff";
            when "10" & x"1b2" => DATA <= x"ffff";
            when "10" & x"1b3" => DATA <= x"ffff";
            when "10" & x"1b4" => DATA <= x"ffff";
            when "10" & x"1b5" => DATA <= x"ffff";
            when "10" & x"1b6" => DATA <= x"ffff";
            when "10" & x"1b7" => DATA <= x"ffff";
            when "10" & x"1b8" => DATA <= x"ffff";
            when "10" & x"1b9" => DATA <= x"ffff";
            when "10" & x"1ba" => DATA <= x"ffff";
            when "10" & x"1bb" => DATA <= x"ffff";
            when "10" & x"1bc" => DATA <= x"ffff";
            when "10" & x"1bd" => DATA <= x"ffff";
            when "10" & x"1be" => DATA <= x"ffff";
            when "10" & x"1bf" => DATA <= x"ffff";
            when "10" & x"1c0" => DATA <= x"ffff";
            when "10" & x"1c1" => DATA <= x"ffff";
            when "10" & x"1c2" => DATA <= x"ffff";
            when "10" & x"1c3" => DATA <= x"ffff";
            when "10" & x"1c4" => DATA <= x"ffff";
            when "10" & x"1c5" => DATA <= x"ffff";
            when "10" & x"1c6" => DATA <= x"ffff";
            when "10" & x"1c7" => DATA <= x"ffff";
            when "10" & x"1c8" => DATA <= x"ffff";
            when "10" & x"1c9" => DATA <= x"ffff";
            when "10" & x"1ca" => DATA <= x"ffff";
            when "10" & x"1cb" => DATA <= x"ffff";
            when "10" & x"1cc" => DATA <= x"ffff";
            when "10" & x"1cd" => DATA <= x"ffff";
            when "10" & x"1ce" => DATA <= x"ffff";
            when "10" & x"1cf" => DATA <= x"ffff";
            when "10" & x"1d0" => DATA <= x"ffff";
            when "10" & x"1d1" => DATA <= x"ffff";
            when "10" & x"1d2" => DATA <= x"ffff";
            when "10" & x"1d3" => DATA <= x"ffff";
            when "10" & x"1d4" => DATA <= x"ffff";
            when "10" & x"1d5" => DATA <= x"ffff";
            when "10" & x"1d6" => DATA <= x"ffff";
            when "10" & x"1d7" => DATA <= x"ffff";
            when "10" & x"1d8" => DATA <= x"ffff";
            when "10" & x"1d9" => DATA <= x"ffff";
            when "10" & x"1da" => DATA <= x"ffff";
            when "10" & x"1db" => DATA <= x"ffff";
            when "10" & x"1dc" => DATA <= x"ffff";
            when "10" & x"1dd" => DATA <= x"ffff";
            when "10" & x"1de" => DATA <= x"ffff";
            when "10" & x"1df" => DATA <= x"ffff";
            when "10" & x"1e0" => DATA <= x"ffff";
            when "10" & x"1e1" => DATA <= x"ffff";
            when "10" & x"1e2" => DATA <= x"ffff";
            when "10" & x"1e3" => DATA <= x"ffff";
            when "10" & x"1e4" => DATA <= x"ffff";
            when "10" & x"1e5" => DATA <= x"ffff";
            when "10" & x"1e6" => DATA <= x"ffff";
            when "10" & x"1e7" => DATA <= x"ffff";
            when "10" & x"1e8" => DATA <= x"ffff";
            when "10" & x"1e9" => DATA <= x"ffff";
            when "10" & x"1ea" => DATA <= x"ffff";
            when "10" & x"1eb" => DATA <= x"ffff";
            when "10" & x"1ec" => DATA <= x"ffff";
            when "10" & x"1ed" => DATA <= x"ffff";
            when "10" & x"1ee" => DATA <= x"ffff";
            when "10" & x"1ef" => DATA <= x"ffff";
            when "10" & x"1f0" => DATA <= x"ffff";
            when "10" & x"1f1" => DATA <= x"ffff";
            when "10" & x"1f2" => DATA <= x"ffff";
            when "10" & x"1f3" => DATA <= x"ffff";
            when "10" & x"1f4" => DATA <= x"ffff";
            when "10" & x"1f5" => DATA <= x"ffff";
            when "10" & x"1f6" => DATA <= x"ffff";
            when "10" & x"1f7" => DATA <= x"ffff";
            when "10" & x"1f8" => DATA <= x"ffff";
            when "10" & x"1f9" => DATA <= x"ffff";
            when "10" & x"1fa" => DATA <= x"ffff";
            when "10" & x"1fb" => DATA <= x"ffff";
            when "10" & x"1fc" => DATA <= x"ffff";
            when "10" & x"1fd" => DATA <= x"ffff";
            when "10" & x"1fe" => DATA <= x"ffff";
            when "10" & x"1ff" => DATA <= x"ffff";
            when "10" & x"200" => DATA <= x"ffff";
            when "10" & x"201" => DATA <= x"ffff";
            when "10" & x"202" => DATA <= x"ffff";
            when "10" & x"203" => DATA <= x"ffff";
            when "10" & x"204" => DATA <= x"ffff";
            when "10" & x"205" => DATA <= x"ffff";
            when "10" & x"206" => DATA <= x"ffff";
            when "10" & x"207" => DATA <= x"ffff";
            when "10" & x"208" => DATA <= x"ffff";
            when "10" & x"209" => DATA <= x"ffff";
            when "10" & x"20a" => DATA <= x"ffff";
            when "10" & x"20b" => DATA <= x"ffff";
            when "10" & x"20c" => DATA <= x"ffff";
            when "10" & x"20d" => DATA <= x"ffff";
            when "10" & x"20e" => DATA <= x"ffff";
            when "10" & x"20f" => DATA <= x"ffff";
            when "10" & x"210" => DATA <= x"ffff";
            when "10" & x"211" => DATA <= x"ffff";
            when "10" & x"212" => DATA <= x"ffff";
            when "10" & x"213" => DATA <= x"ffff";
            when "10" & x"214" => DATA <= x"ffff";
            when "10" & x"215" => DATA <= x"ffff";
            when "10" & x"216" => DATA <= x"ffff";
            when "10" & x"217" => DATA <= x"ffff";
            when "10" & x"218" => DATA <= x"ffff";
            when "10" & x"219" => DATA <= x"ffff";
            when "10" & x"21a" => DATA <= x"ffff";
            when "10" & x"21b" => DATA <= x"ffff";
            when "10" & x"21c" => DATA <= x"ffff";
            when "10" & x"21d" => DATA <= x"ffff";
            when "10" & x"21e" => DATA <= x"ffff";
            when "10" & x"21f" => DATA <= x"ffff";
            when "10" & x"220" => DATA <= x"ffff";
            when "10" & x"221" => DATA <= x"ffff";
            when "10" & x"222" => DATA <= x"ffff";
            when "10" & x"223" => DATA <= x"ffff";
            when "10" & x"224" => DATA <= x"ffff";
            when "10" & x"225" => DATA <= x"ffff";
            when "10" & x"226" => DATA <= x"ffff";
            when "10" & x"227" => DATA <= x"ffff";
            when "10" & x"228" => DATA <= x"ffff";
            when "10" & x"229" => DATA <= x"ffff";
            when "10" & x"22a" => DATA <= x"ffff";
            when "10" & x"22b" => DATA <= x"ffff";
            when "10" & x"22c" => DATA <= x"ffff";
            when "10" & x"22d" => DATA <= x"ffff";
            when "10" & x"22e" => DATA <= x"ffff";
            when "10" & x"22f" => DATA <= x"ffff";
            when "10" & x"230" => DATA <= x"ffff";
            when "10" & x"231" => DATA <= x"ffff";
            when "10" & x"232" => DATA <= x"ffff";
            when "10" & x"233" => DATA <= x"ffff";
            when "10" & x"234" => DATA <= x"ffff";
            when "10" & x"235" => DATA <= x"ffff";
            when "10" & x"236" => DATA <= x"ffff";
            when "10" & x"237" => DATA <= x"ffff";
            when "10" & x"238" => DATA <= x"ffff";
            when "10" & x"239" => DATA <= x"ffff";
            when "10" & x"23a" => DATA <= x"ffff";
            when "10" & x"23b" => DATA <= x"ffff";
            when "10" & x"23c" => DATA <= x"ffff";
            when "10" & x"23d" => DATA <= x"ffff";
            when "10" & x"23e" => DATA <= x"ffff";
            when "10" & x"23f" => DATA <= x"ffff";
            when "10" & x"240" => DATA <= x"ffff";
            when "10" & x"241" => DATA <= x"ffff";
            when "10" & x"242" => DATA <= x"ffff";
            when "10" & x"243" => DATA <= x"ffff";
            when "10" & x"244" => DATA <= x"ffff";
            when "10" & x"245" => DATA <= x"ffff";
            when "10" & x"246" => DATA <= x"ffff";
            when "10" & x"247" => DATA <= x"ffff";
            when "10" & x"248" => DATA <= x"ffff";
            when "10" & x"249" => DATA <= x"ffff";
            when "10" & x"24a" => DATA <= x"ffff";
            when "10" & x"24b" => DATA <= x"ffff";
            when "10" & x"24c" => DATA <= x"ffff";
            when "10" & x"24d" => DATA <= x"ffff";
            when "10" & x"24e" => DATA <= x"ffff";
            when "10" & x"24f" => DATA <= x"ffff";
            when "10" & x"250" => DATA <= x"ffff";
            when "10" & x"251" => DATA <= x"1000";
            when "10" & x"252" => DATA <= x"e0e0";
            when "10" & x"253" => DATA <= x"e0e0";
            when "10" & x"254" => DATA <= x"e0e0";
            when "10" & x"255" => DATA <= x"e0e0";
            when "10" & x"256" => DATA <= x"80c0";
            when "10" & x"257" => DATA <= x"0004";
            when "10" & x"258" => DATA <= x"2400";
            when "10" & x"259" => DATA <= x"081e";
            when "10" & x"25a" => DATA <= x"a00a";
            when "10" & x"25b" => DATA <= x"ff74";
            when "10" & x"25c" => DATA <= x"5000";
            when "10" & x"25d" => DATA <= x"3e80";
            when "10" & x"25e" => DATA <= x"1fe0";
            when "10" & x"25f" => DATA <= x"6aff";
            when "10" & x"260" => DATA <= x"7c20";
            when "10" & x"261" => DATA <= x"2801";
            when "10" & x"262" => DATA <= x"fe00";
            when "10" & x"263" => DATA <= x"6f8b";
            when "10" & x"264" => DATA <= x"ebfe";
            when "10" & x"265" => DATA <= x"801f";
            when "10" & x"266" => DATA <= x"ec00";
            when "10" & x"267" => DATA <= x"f980";
            when "10" & x"268" => DATA <= x"1e3f";
            when "10" & x"269" => DATA <= x"a007";
            when "10" & x"26a" => DATA <= x"fb6d";
            when "10" & x"26b" => DATA <= x"fce0";
            when "10" & x"26c" => DATA <= x"9007";
            when "10" & x"26d" => DATA <= x"f802";
            when "10" & x"26e" => DATA <= x"bfeb";
            when "10" & x"26f" => DATA <= x"e280";
            when "10" & x"270" => DATA <= x"1fe0";
            when "10" & x"271" => DATA <= x"07f8";
            when "10" & x"272" => DATA <= x"1cbe";
            when "10" & x"273" => DATA <= x"ffa0";
            when "10" & x"274" => DATA <= x"07fb";
            when "10" & x"275" => DATA <= x"81fe";
            when "10" & x"276" => DATA <= x"ac00";
            when "10" & x"277" => DATA <= x"27e8";
            when "10" & x"278" => DATA <= x"03bf";
            when "10" & x"279" => DATA <= x"de35";
            when "10" & x"27a" => DATA <= x"8140";
            when "10" & x"27b" => DATA <= x"17ff";
            when "10" & x"27c" => DATA <= x"400f";
            when "10" & x"27d" => DATA <= x"f014";
            when "10" & x"27e" => DATA <= x"ffd0";
            when "10" & x"27f" => DATA <= x"03fd";
            when "10" & x"280" => DATA <= x"e0ff";
            when "10" & x"281" => DATA <= x"7800";
            when "10" & x"282" => DATA <= x"c1f4";
            when "10" & x"283" => DATA <= x"00ff";
            when "10" & x"284" => DATA <= x"00bf";
            when "10" & x"285" => DATA <= x"d408";
            when "10" & x"286" => DATA <= x"071d";
            when "10" & x"287" => DATA <= x"005f";
            when "10" & x"288" => DATA <= x"fd00";
            when "10" & x"289" => DATA <= x"3fd7";
            when "10" & x"28a" => DATA <= x"f3ff";
            when "10" & x"28b" => DATA <= x"400f";
            when "10" & x"28c" => DATA <= x"f7d4";
            when "10" & x"28d" => DATA <= x"ffd0";
            when "10" & x"28e" => DATA <= x"03fc";
            when "10" & x"28f" => DATA <= x"00ff";
            when "10" & x"290" => DATA <= x"080c";
            when "10" & x"291" => DATA <= x"c474";
            when "10" & x"292" => DATA <= x"00ff";
            when "10" & x"293" => DATA <= x"403f";
            when "10" & x"294" => DATA <= x"df8f";
            when "10" & x"295" => DATA <= x"f7f5";
            when "10" & x"296" => DATA <= x"003f";
            when "10" & x"297" => DATA <= x"dfd3";
            when "10" & x"298" => DATA <= x"ff40";
            when "10" & x"299" => DATA <= x"0ff7";
            when "10" & x"29a" => DATA <= x"ecff";
            when "10" & x"29b" => DATA <= x"d003";
            when "10" & x"29c" => DATA <= x"fc00";
            when "10" & x"29d" => DATA <= x"ff20";
            when "10" & x"29e" => DATA <= x"bbd9";
            when "10" & x"29f" => DATA <= x"f400";
            when "10" & x"2a0" => DATA <= x"ff00";
            when "10" & x"2a1" => DATA <= x"3fde";
            when "10" & x"2a2" => DATA <= x"0fe7";
            when "10" & x"2a3" => DATA <= x"e500";
            when "10" & x"2a4" => DATA <= x"5ffd";
            when "10" & x"2a5" => DATA <= x"003f";
            when "10" & x"2a6" => DATA <= x"cff3";
            when "10" & x"2a7" => DATA <= x"ff40";
            when "10" & x"2a8" => DATA <= x"0ff0";
            when "10" & x"2a9" => DATA <= x"03fc";
            when "10" & x"2aa" => DATA <= x"82e7";
            when "10" & x"2ab" => DATA <= x"23d0";
            when "10" & x"2ac" => DATA <= x"03fc";
            when "10" & x"2ad" => DATA <= x"00ff";
            when "10" & x"2ae" => DATA <= x"7057";
            when "10" & x"2af" => DATA <= x"e500";
            when "10" & x"2b0" => DATA <= x"3fdf";
            when "10" & x"2b1" => DATA <= x"13ff";
            when "10" & x"2b2" => DATA <= x"4017";
            when "10" & x"2b3" => DATA <= x"ff40";
            when "10" & x"2b4" => DATA <= x"0ff0";
            when "10" & x"2b5" => DATA <= x"3bfc";
            when "10" & x"2b6" => DATA <= x"7eff";
            when "10" & x"2b7" => DATA <= x"3fd0";
            when "10" & x"2b8" => DATA <= x"03fc";
            when "10" & x"2b9" => DATA <= x"00ff";
            when "10" & x"2ba" => DATA <= x"0033";
            when "10" & x"2bb" => DATA <= x"9814";
            when "10" & x"2bc" => DATA <= x"00ff";
            when "10" & x"2bd" => DATA <= x"003f";
            when "10" & x"2be" => DATA <= x"df95";
            when "10" & x"2bf" => DATA <= x"ff40";
            when "10" & x"2c0" => DATA <= x"0ff7";
            when "10" & x"2c1" => DATA <= x"f4ff";
            when "10" & x"2c2" => DATA <= x"d005";
            when "10" & x"2c3" => DATA <= x"ffd0";
            when "10" & x"2c4" => DATA <= x"05ff";
            when "10" & x"2c5" => DATA <= x"d005";
            when "10" & x"2c6" => DATA <= x"ffd0";
            when "10" & x"2c7" => DATA <= x"05ff";
            when "10" & x"2c8" => DATA <= x"d005";
            when "10" & x"2c9" => DATA <= x"ffd0";
            when "10" & x"2ca" => DATA <= x"077f";
            when "10" & x"2cb" => DATA <= x"d3f8";
            when "10" & x"2cc" => DATA <= x"fe80";
            when "10" & x"2cd" => DATA <= x"27fd";
            when "10" & x"2ce" => DATA <= x"9ce0";
            when "10" & x"2cf" => DATA <= x"a00b";
            when "10" & x"2d0" => DATA <= x"ffa0";
            when "10" & x"2d1" => DATA <= x"0eff";
            when "10" & x"2d2" => DATA <= x"3fa7";
            when "10" & x"2d3" => DATA <= x"c1f4";
            when "10" & x"2d4" => DATA <= x"013f";
            when "10" & x"2d5" => DATA <= x"efb7";
            when "10" & x"2d6" => DATA <= x"cd00";
            when "10" & x"2d7" => DATA <= x"6ff9";
            when "10" & x"2d8" => DATA <= x"7e80";
            when "10" & x"2d9" => DATA <= x"37fd";
            when "10" & x"2da" => DATA <= x"ed40";
            when "10" & x"2db" => DATA <= x"1bfe";
            when "10" & x"2dc" => DATA <= x"17a0";
            when "10" & x"2dd" => DATA <= x"0dff";
            when "10" & x"2de" => DATA <= x"7ed0";
            when "10" & x"2df" => DATA <= x"06ff";
            when "10" & x"2e0" => DATA <= x"9fe8";
            when "10" & x"2e1" => DATA <= x"037f";
            when "10" & x"2e2" => DATA <= x"f803";
            when "10" & x"2e3" => DATA <= x"bfdf";
            when "10" & x"2e4" => DATA <= x"ad84";
            when "10" & x"2e5" => DATA <= x"0500";
            when "10" & x"2e6" => DATA <= x"4ffb";
            when "10" & x"2e7" => DATA <= x"01bb";
            when "10" & x"2e8" => DATA <= x"400f";
            when "10" & x"2e9" => DATA <= x"f3fc";
            when "10" & x"2ea" => DATA <= x"ffd0";
            when "10" & x"2eb" => DATA <= x"03fc";
            when "10" & x"2ec" => DATA <= x"ffdf";
            when "10" & x"2ed" => DATA <= x"e2fa";
            when "10" & x"2ee" => DATA <= x"007f";
            when "10" & x"2ef" => DATA <= x"801f";
            when "10" & x"2f0" => DATA <= x"e417";
            when "10" & x"2f1" => DATA <= x"3f00";
            when "10" & x"2f2" => DATA <= x"3fc0";
            when "10" & x"2f3" => DATA <= x"0ff6";
            when "10" & x"2f4" => DATA <= x"03f9";
            when "10" & x"2f5" => DATA <= x"f140";
            when "10" & x"2f6" => DATA <= x"17ff";
            when "10" & x"2f7" => DATA <= x"400f";
            when "10" & x"2f8" => DATA <= x"f6fc";
            when "10" & x"2f9" => DATA <= x"ffd0";
            when "10" & x"2fa" => DATA <= x"03fc";
            when "10" & x"2fb" => DATA <= x"3fdf";
            when "10" & x"2fc" => DATA <= x"e7fa";
            when "10" & x"2fd" => DATA <= x"007f";
            when "10" & x"2fe" => DATA <= x"a01f";
            when "10" & x"2ff" => DATA <= x"e876";
            when "10" & x"300" => DATA <= x"ff00";
            when "10" & x"301" => DATA <= x"3fc0";
            when "10" & x"302" => DATA <= x"eff7";
            when "10" & x"303" => DATA <= x"5bfd";
            when "10" & x"304" => DATA <= x"c140";
            when "10" & x"305" => DATA <= x"0ff7";
            when "10" & x"306" => DATA <= x"44ff";
            when "10" & x"307" => DATA <= x"d003";
            when "10" & x"308" => DATA <= x"fc00";
            when "10" & x"309" => DATA <= x"ff1f";
            when "10" & x"30a" => DATA <= x"bfc7";
            when "10" & x"30b" => DATA <= x"f400";
            when "10" & x"30c" => DATA <= x"ff40";
            when "10" & x"30d" => DATA <= x"3fc9";
            when "10" & x"30e" => DATA <= x"0ec7";
            when "10" & x"30f" => DATA <= x"2500";
            when "10" & x"310" => DATA <= x"3fc0";
            when "10" & x"311" => DATA <= x"f3ff";
            when "10" & x"312" => DATA <= x"400f";
            when "10" & x"313" => DATA <= x"f5ac";
            when "10" & x"314" => DATA <= x"ffd0";
            when "10" & x"315" => DATA <= x"03fc";
            when "10" & x"316" => DATA <= x"02ff";
            when "10" & x"317" => DATA <= x"03b7";
            when "10" & x"318" => DATA <= x"cc74";
            when "10" & x"319" => DATA <= x"00ff";
            when "10" & x"31a" => DATA <= x"603f";
            when "10" & x"31b" => DATA <= x"d82f";
            when "10" & x"31c" => DATA <= x"f6e5";
            when "10" & x"31d" => DATA <= x"003f";
            when "10" & x"31e" => DATA <= x"c06f";
            when "10" & x"31f" => DATA <= x"f7dd";
            when "10" & x"320" => DATA <= x"7fd0";
            when "10" & x"321" => DATA <= x"03fd";
            when "10" & x"322" => DATA <= x"f93f";
            when "10" & x"323" => DATA <= x"f400";
            when "10" & x"324" => DATA <= x"ff1f";
            when "10" & x"325" => DATA <= x"bfe8";
            when "10" & x"326" => DATA <= x"3c0f";
            when "10" & x"327" => DATA <= x"400f";
            when "10" & x"328" => DATA <= x"f503";
            when "10" & x"329" => DATA <= x"fd10";
            when "10" & x"32a" => DATA <= x"d778";
            when "10" & x"32b" => DATA <= x"5003";
            when "10" & x"32c" => DATA <= x"fc06";
            when "10" & x"32d" => DATA <= x"ff7d";
            when "10" & x"32e" => DATA <= x"d7fd";
            when "10" & x"32f" => DATA <= x"003f";
            when "10" & x"330" => DATA <= x"dc13";
            when "10" & x"331" => DATA <= x"ff40";
            when "10" & x"332" => DATA <= x"0ff1";
            when "10" & x"333" => DATA <= x"fbfc";
            when "10" & x"334" => DATA <= x"1e07";
            when "10" & x"335" => DATA <= x"e007";
            when "10" & x"336" => DATA <= x"f8c1";
            when "10" & x"337" => DATA <= x"8610";
            when "10" & x"338" => DATA <= x"00bc";
            when "10" & x"339" => DATA <= x"2801";
            when "10" & x"33a" => DATA <= x"fe00";
            when "10" & x"33b" => DATA <= x"78bc";
            when "10" & x"33c" => DATA <= x"2bfe";
            when "10" & x"33d" => DATA <= x"801f";
            when "10" & x"33e" => DATA <= x"af0e";
            when "10" & x"33f" => DATA <= x"ff3f";
            when "10" & x"340" => DATA <= x"d007";
            when "10" & x"341" => DATA <= x"7f97";
            when "10" & x"342" => DATA <= x"c07c";
            when "10" & x"343" => DATA <= x"00ff";
            when "10" & x"344" => DATA <= x"1fa0";
            when "10" & x"345" => DATA <= x"c20c";
            when "10" & x"346" => DATA <= x"07a5";
            when "10" & x"347" => DATA <= x"0000";
            when "10" & x"348" => DATA <= x"4000";
            when "10" & x"349" => DATA <= x"1205";
            when "10" & x"34a" => DATA <= x"3887";
            when "10" & x"34b" => DATA <= x"8381";
            when "10" & x"34c" => DATA <= x"e0e0";
            when "10" & x"34d" => DATA <= x"7839";
            when "10" & x"34e" => DATA <= x"43db";
            when "10" & x"34f" => DATA <= x"df5f";
            when "10" & x"350" => DATA <= x"eef0";
            when "10" & x"351" => DATA <= x"051f";
            when "10" & x"352" => DATA <= x"0fc7";
            when "10" & x"353" => DATA <= x"d47e";
            when "10" & x"354" => DATA <= x"3e78";
            when "10" & x"355" => DATA <= x"3000";
            when "10" & x"356" => DATA <= x"0181";
            when "10" & x"357" => DATA <= x"c57c";
            when "10" & x"358" => DATA <= x"5000";
            when "10" & x"359" => DATA <= x"0dfc";
            when "10" & x"35a" => DATA <= x"f060";
            when "10" & x"35b" => DATA <= x"20df";
            when "10" & x"35c" => DATA <= x"f401";
            when "10" & x"35d" => DATA <= x"c61d";
            when "10" & x"35e" => DATA <= x"6090";
            when "10" & x"35f" => DATA <= x"6020";
            when "10" & x"360" => DATA <= x"0003";
            when "10" & x"361" => DATA <= x"0385";
            when "10" & x"362" => DATA <= x"7800";
            when "10" & x"363" => DATA <= x"0020";
            when "10" & x"364" => DATA <= x"77e3";
            when "10" & x"365" => DATA <= x"8100";
            when "10" & x"366" => DATA <= x"8107";
            when "10" & x"367" => DATA <= x"8008";
            when "10" & x"368" => DATA <= x"0607";
            when "10" & x"369" => DATA <= x"0cb0";
            when "10" & x"36a" => DATA <= x"8838";
            when "10" & x"36b" => DATA <= x"00c1";
            when "10" & x"36c" => DATA <= x"dc00";
            when "10" & x"36d" => DATA <= x"0010";
            when "10" & x"36e" => DATA <= x"39f0";
            when "10" & x"36f" => DATA <= x"c040";
            when "10" & x"370" => DATA <= x"00c1";
            when "10" & x"371" => DATA <= x"e00a";
            when "10" & x"372" => DATA <= x"c09c";
            when "10" & x"373" => DATA <= x"341f";
            when "10" & x"374" => DATA <= x"0030";
            when "10" & x"375" => DATA <= x"502c";
            when "10" & x"376" => DATA <= x"0403";
            when "10" & x"377" => DATA <= x"0380";
            when "10" & x"378" => DATA <= x"1820";
            when "10" & x"379" => DATA <= x"3038";
            when "10" & x"37a" => DATA <= x"3c7f";
            when "10" & x"37b" => DATA <= x"c014";
            when "10" & x"37c" => DATA <= x"1e0e";
            when "10" & x"37d" => DATA <= x"a0c0";
            when "10" & x"37e" => DATA <= x"073f";
            when "10" & x"37f" => DATA <= x"90f8";
            when "10" & x"380" => DATA <= x"4c22";
            when "10" & x"381" => DATA <= x"f500";
            when "10" & x"382" => DATA <= x"5080";
            when "10" & x"383" => DATA <= x"02b8";
            when "10" & x"384" => DATA <= x"1e00";
            when "10" & x"385" => DATA <= x"7000";
            when "10" & x"386" => DATA <= x"7c1e";
            when "10" & x"387" => DATA <= x"1f1f";
            when "10" & x"388" => DATA <= x"9fc3";
            when "10" & x"389" => DATA <= x"fdfc";
            when "10" & x"38a" => DATA <= x"fca3";
            when "10" & x"38b" => DATA <= x"81e0";
            when "10" & x"38c" => DATA <= x"01fe";
            when "10" & x"38d" => DATA <= x"2b41";
            when "10" & x"38e" => DATA <= x"80fa";
            when "10" & x"38f" => DATA <= x"0004";
            when "10" & x"390" => DATA <= x"ff50";
            when "10" & x"391" => DATA <= x"0428";
            when "10" & x"392" => DATA <= x"0021";
            when "10" & x"393" => DATA <= x"4000";
            when "10" & x"394" => DATA <= x"707f";
            when "10" & x"395" => DATA <= x"0f87";
            when "10" & x"396" => DATA <= x"87e8";
            when "10" & x"397" => DATA <= x"07e0";
            when "10" & x"398" => DATA <= x"028f";
            when "10" & x"399" => DATA <= x"28e0";
            when "10" & x"39a" => DATA <= x"78ff";
            when "10" & x"39b" => DATA <= x"7ef6";
            when "10" & x"39c" => DATA <= x"0309";
            when "10" & x"39d" => DATA <= x"00c0";
            when "10" & x"39e" => DATA <= x"21d0";
            when "10" & x"39f" => DATA <= x"0ef0";
            when "10" & x"3a0" => DATA <= x"8068";
            when "10" & x"3a1" => DATA <= x"000e";
            when "10" & x"3a2" => DATA <= x"83a8";
            when "10" & x"3a3" => DATA <= x"1618";
            when "10" & x"3a4" => DATA <= x"0180";
            when "10" & x"3a5" => DATA <= x"c163";
            when "10" & x"3a6" => DATA <= x"d43a";
            when "10" & x"3a7" => DATA <= x"7dfe";
            when "10" & x"3a8" => DATA <= x"00ef";
            when "10" & x"3a9" => DATA <= x"f5a5";
            when "10" & x"3aa" => DATA <= x"4a00";
            when "10" & x"3ab" => DATA <= x"0edc";
            when "10" & x"3ac" => DATA <= x"1e07";
            when "10" & x"3ad" => DATA <= x"0257";
            when "10" & x"3ae" => DATA <= x"2804";
            when "10" & x"3af" => DATA <= x"3c3e";
            when "10" & x"3b0" => DATA <= x"1f87";
            when "10" & x"3b1" => DATA <= x"f83f";
            when "10" & x"3b2" => DATA <= x"8038";
            when "10" & x"3b3" => DATA <= x"603c";
            when "10" & x"3b4" => DATA <= x"1f00";
            when "10" & x"3b5" => DATA <= x"7830";
            when "10" & x"3b6" => DATA <= x"0820";
            when "10" & x"3b7" => DATA <= x"7eaf";
            when "10" & x"3b8" => DATA <= x"e3f5";
            when "10" & x"3b9" => DATA <= x"7f70";
            when "10" & x"3ba" => DATA <= x"057f";
            when "10" & x"3bb" => DATA <= x"f1f8";
            when "10" & x"3bc" => DATA <= x"02bf";
            when "10" & x"3bd" => DATA <= x"1faf";
            when "10" & x"3be" => DATA <= x"f005";
            when "10" & x"3bf" => DATA <= x"0400";
            when "10" & x"3c0" => DATA <= x"2bfd";
            when "10" & x"3c1" => DATA <= x"ee37";
            when "10" & x"3c2" => DATA <= x"1408";
            when "10" & x"3c3" => DATA <= x"4041";
            when "10" & x"3c4" => DATA <= x"0aff";
            when "10" & x"3c5" => DATA <= x"7f00";
            when "10" & x"3c6" => DATA <= x"40a9";
            when "10" & x"3c7" => DATA <= x"9038";
            when "10" & x"3c8" => DATA <= x"21fe";
            when "10" & x"3c9" => DATA <= x"3f0f";
            when "10" & x"3ca" => DATA <= x"f008";
            when "10" & x"3cb" => DATA <= x"1444";
            when "10" & x"3cc" => DATA <= x"3fa3";
            when "10" & x"3cd" => DATA <= x"e0f0";
            when "10" & x"3ce" => DATA <= x"3a83";
            when "10" & x"3cf" => DATA <= x"000e";
            when "10" & x"3d0" => DATA <= x"0381";
            when "10" & x"3d1" => DATA <= x"e1f8";
            when "10" & x"3d2" => DATA <= x"f87e";
            when "10" & x"3d3" => DATA <= x"1f80";
            when "10" & x"3d4" => DATA <= x"0ffa";
            when "10" & x"3d5" => DATA <= x"00ef";
            when "10" & x"3d6" => DATA <= x"fa00";
            when "10" & x"3d7" => DATA <= x"e1f0";
            when "10" & x"3d8" => DATA <= x"7f03";
            when "10" & x"3d9" => DATA <= x"801e";
            when "10" & x"3da" => DATA <= x"0180";
            when "10" & x"3db" => DATA <= x"e70f";
            when "10" & x"3dc" => DATA <= x"07c0";
            when "10" & x"3dd" => DATA <= x"07fb";
            when "10" & x"3de" => DATA <= x"0030";
            when "10" & x"3df" => DATA <= x"2da8";
            when "10" & x"3e0" => DATA <= x"c340";
            when "10" & x"3e1" => DATA <= x"02b4";
            when "10" & x"3e2" => DATA <= x"0806";
            when "10" & x"3e3" => DATA <= x"9007";
            when "10" & x"3e4" => DATA <= x"ef00";
            when "10" & x"3e5" => DATA <= x"0400";
            when "10" & x"3e6" => DATA <= x"9400";
            when "10" & x"3e7" => DATA <= x"bfb0";
            when "10" & x"3e8" => DATA <= x"0008";
            when "10" & x"3e9" => DATA <= x"fde0";
            when "10" & x"3ea" => DATA <= x"f83c";
            when "10" & x"3eb" => DATA <= x"71c7";
            when "10" & x"3ec" => DATA <= x"0077";
            when "10" & x"3ed" => DATA <= x"03c1";
            when "10" & x"3ee" => DATA <= x"f200";
            when "10" & x"3ef" => DATA <= x"2058";
            when "10" & x"3f0" => DATA <= x"8001";
            when "10" & x"3f1" => DATA <= x"faf8";
            when "10" & x"3f2" => DATA <= x"4870";
            when "10" & x"3f3" => DATA <= x"0004";
            when "10" & x"3f4" => DATA <= x"00f7";
            when "10" & x"3f5" => DATA <= x"0057";
            when "10" & x"3f6" => DATA <= x"8538";
            when "10" & x"3f7" => DATA <= x"0c0e";
            when "10" & x"3f8" => DATA <= x"1406";
            when "10" & x"3f9" => DATA <= x"c160";
            when "10" & x"3fa" => DATA <= x"5703";
            when "10" & x"3fb" => DATA <= x"e5f8";
            when "10" & x"3fc" => DATA <= x"fa70";
            when "10" & x"3fd" => DATA <= x"5f1b";
            when "10" & x"3fe" => DATA <= x"ff7c";
            when "10" & x"3ff" => DATA <= x"deef";
            when "10" & x"400" => DATA <= x"37ff";
            when "10" & x"401" => DATA <= x"bfb7";
            when "10" & x"402" => DATA <= x"c013";
            when "10" & x"403" => DATA <= x"0150";
            when "10" & x"404" => DATA <= x"4070";
            when "10" & x"405" => DATA <= x"407c";
            when "10" & x"406" => DATA <= x"1f40";
            when "10" & x"407" => DATA <= x"e0f5";
            when "10" & x"408" => DATA <= x"fb20";
            when "10" & x"409" => DATA <= x"0141";
            when "10" & x"40a" => DATA <= x"c0c0";
            when "10" & x"40b" => DATA <= x"7707";
            when "10" & x"40c" => DATA <= x"f800";
            when "10" & x"40d" => DATA <= x"4060";
            when "10" & x"40e" => DATA <= x"3f0f";
            when "10" & x"40f" => DATA <= x"d07a";
            when "10" & x"410" => DATA <= x"1f80";
            when "10" & x"411" => DATA <= x"0314";
            when "10" & x"412" => DATA <= x"381e";
            when "10" & x"413" => DATA <= x"0f80";
            when "10" & x"414" => DATA <= x"3c18";
            when "10" & x"415" => DATA <= x"04a0";
            when "10" & x"416" => DATA <= x"703f";
            when "10" & x"417" => DATA <= x"87c1";
            when "10" & x"418" => DATA <= x"e070";
            when "10" & x"419" => DATA <= x"1a80";
            when "10" & x"41a" => DATA <= x"0022";
            when "10" & x"41b" => DATA <= x"0380";
            when "10" & x"41c" => DATA <= x"e078";
            when "10" & x"41d" => DATA <= x"3f00";
            when "10" & x"41e" => DATA <= x"2228";
            when "10" & x"41f" => DATA <= x"6018";
            when "10" & x"420" => DATA <= x"1c04";
            when "10" & x"421" => DATA <= x"0602";
            when "10" & x"422" => DATA <= x"0fd0";
            when "10" & x"423" => DATA <= x"1389";
            when "10" & x"424" => DATA <= x"c0e2";
            when "10" & x"425" => DATA <= x"7038";
            when "10" & x"426" => DATA <= x"9fcf";
            when "10" & x"427" => DATA <= x"f3c0";
            when "10" & x"428" => DATA <= x"fc0e";
            when "10" & x"429" => DATA <= x"0140";
            when "10" & x"42a" => DATA <= x"b801";
            when "10" & x"42b" => DATA <= x"a01a";
            when "10" & x"42c" => DATA <= x"0003";
            when "10" & x"42d" => DATA <= x"01c8";
            when "10" & x"42e" => DATA <= x"e070";
            when "10" & x"42f" => DATA <= x"0010";
            when "10" & x"430" => DATA <= x"0084";
            when "10" & x"431" => DATA <= x"a804";
            when "10" & x"432" => DATA <= x"2200";
            when "10" & x"433" => DATA <= x"000f";
            when "10" & x"434" => DATA <= x"1fbf";
            when "10" & x"435" => DATA <= x"c3e0";
            when "10" & x"436" => DATA <= x"701b";
            when "10" & x"437" => DATA <= x"8640";
            when "10" & x"438" => DATA <= x"0100";
            when "10" & x"439" => DATA <= x"ca0f";
            when "10" & x"43a" => DATA <= x"e004";
            when "10" & x"43b" => DATA <= x"1d01";
            when "10" & x"43c" => DATA <= x"a0c0";
            when "10" & x"43d" => DATA <= x"601a";
            when "10" & x"43e" => DATA <= x"ffaf";
            when "10" & x"43f" => DATA <= x"81c0";
            when "10" & x"440" => DATA <= x"6110";
            when "10" & x"441" => DATA <= x"007f";
            when "10" & x"442" => DATA <= x"80c1";
            when "10" & x"443" => DATA <= x"e006";
            when "10" & x"444" => DATA <= x"03c1";
            when "10" & x"445" => DATA <= x"fefe";
            when "10" & x"446" => DATA <= x"03d0";
            when "10" & x"447" => DATA <= x"0480";
            when "10" & x"448" => DATA <= x"9fd8";
            when "10" & x"449" => DATA <= x"0de9";
            when "10" & x"44a" => DATA <= x"dfaf";
            when "10" & x"44b" => DATA <= x"fbf7";
            when "10" & x"44c" => DATA <= x"afff";
            when "10" & x"44d" => DATA <= x"7138";
            when "10" & x"44e" => DATA <= x"87a8";
            when "10" & x"44f" => DATA <= x"703c";
            when "10" & x"450" => DATA <= x"1ca0";
            when "10" & x"451" => DATA <= x"0026";
            when "10" & x"452" => DATA <= x"f7bb";
            when "10" & x"453" => DATA <= x"8000";
            when "10" & x"454" => DATA <= x"74f5";
            when "10" & x"455" => DATA <= x"5d2f";
            when "10" & x"456" => DATA <= x"9fc1";
            when "10" & x"457" => DATA <= x"ea00";
            when "10" & x"458" => DATA <= x"2857";
            when "10" & x"459" => DATA <= x"fbed";
            when "10" & x"45a" => DATA <= x"fe00";
            when "10" & x"45b" => DATA <= x"7e50";
            when "10" & x"45c" => DATA <= x"02fc";
            when "10" & x"45d" => DATA <= x"fcff";
            when "10" & x"45e" => DATA <= x"6780";
            when "10" & x"45f" => DATA <= x"0fef";
            when "10" & x"460" => DATA <= x"f48f";
            when "10" & x"461" => DATA <= x"7fbd";
            when "10" & x"462" => DATA <= x"1e0e";
            when "10" & x"463" => DATA <= x"0780";
            when "10" & x"464" => DATA <= x"03bf";
            when "10" & x"465" => DATA <= x"c7e7";
            when "10" & x"466" => DATA <= x"f3e8";
            when "10" & x"467" => DATA <= x"fc04";
            when "10" & x"468" => DATA <= x"ff7e";
            when "10" & x"469" => DATA <= x"bfd0";
            when "10" & x"46a" => DATA <= x"8637";
            when "10" & x"46b" => DATA <= x"9a40";
            when "10" & x"46c" => DATA <= x"415f";
            when "10" & x"46d" => DATA <= x"d47e";
            when "10" & x"46e" => DATA <= x"0203";
            when "10" & x"46f" => DATA <= x"a218";
            when "10" & x"470" => DATA <= x"35fe";
            when "10" & x"471" => DATA <= x"fe4f";
            when "10" & x"472" => DATA <= x"1000";
            when "10" & x"473" => DATA <= x"0040";
            when "10" & x"474" => DATA <= x"2afd";
            when "10" & x"475" => DATA <= x"feef";
            when "10" & x"476" => DATA <= x"1d80";
            when "10" & x"477" => DATA <= x"a800";
            when "10" & x"478" => DATA <= x"c15f";
            when "10" & x"479" => DATA <= x"aff7";
            when "10" & x"47a" => DATA <= x"f235";
            when "10" & x"47b" => DATA <= x"98c4";
            when "10" & x"47c" => DATA <= x"0157";
            when "10" & x"47d" => DATA <= x"fafd";
            when "10" & x"47e" => DATA <= x"fe14";
            when "10" & x"47f" => DATA <= x"0008";
            when "10" & x"480" => DATA <= x"0167";
            when "10" & x"481" => DATA <= x"f77a";
            when "10" & x"482" => DATA <= x"fc66";
            when "10" & x"483" => DATA <= x"0024";
            when "10" & x"484" => DATA <= x"1018";
            when "10" & x"485" => DATA <= x"0fb7";
            when "10" & x"486" => DATA <= x"bbfd";
            when "10" & x"487" => DATA <= x"f800";
            when "10" & x"488" => DATA <= x"45b2";
            when "10" & x"489" => DATA <= x"c21d";
            when "10" & x"48a" => DATA <= x"fe8f";
            when "10" & x"48b" => DATA <= x"4000";
            when "10" & x"48c" => DATA <= x"1000";
            when "10" & x"48d" => DATA <= x"077d";
            when "10" & x"48e" => DATA <= x"7fa9";
            when "10" & x"48f" => DATA <= x"c0e0";
            when "10" & x"490" => DATA <= x"0020";
            when "10" & x"491" => DATA <= x"03bf";
            when "10" & x"492" => DATA <= x"dee0";
            when "10" & x"493" => DATA <= x"4000";
            when "10" & x"494" => DATA <= x"9009";
            when "10" & x"495" => DATA <= x"3fe0";
            when "10" & x"496" => DATA <= x"0641";
            when "10" & x"497" => DATA <= x"0d00";
            when "10" & x"498" => DATA <= x"ff77";
            when "10" & x"499" => DATA <= x"bfcf";
            when "10" & x"49a" => DATA <= x"e000";
            when "10" & x"49b" => DATA <= x"1098";
            when "10" & x"49c" => DATA <= x"00ef";
            when "10" & x"49d" => DATA <= x"aff7";
            when "10" & x"49e" => DATA <= x"0000";
            when "10" & x"49f" => DATA <= x"0844";
            when "10" & x"4a0" => DATA <= x"003f";
            when "10" & x"4a1" => DATA <= x"5eaf";
            when "10" & x"4a2" => DATA <= x"d7fb";
            when "10" & x"4a3" => DATA <= x"0000";
            when "10" & x"4a4" => DATA <= x"0a02";
            when "10" & x"4a5" => DATA <= x"77fb";
            when "10" & x"4a6" => DATA <= x"e480";
            when "10" & x"4a7" => DATA <= x"0700";
            when "10" & x"4a8" => DATA <= x"007b";
            when "10" & x"4a9" => DATA <= x"fd02";
            when "10" & x"4aa" => DATA <= x"4800";
            when "10" & x"4ab" => DATA <= x"1202";
            when "10" & x"4ac" => DATA <= x"6bf6";
            when "10" & x"4ad" => DATA <= x"fbfc";
            when "10" & x"4ae" => DATA <= x"661a";
            when "10" & x"4af" => DATA <= x"a007";
            when "10" & x"4b0" => DATA <= x"03f5";
            when "10" & x"4b1" => DATA <= x"deff";
            when "10" & x"4b2" => DATA <= x"7d00";
            when "10" & x"4b3" => DATA <= x"0482";
            when "10" & x"4b4" => DATA <= x"1211";
            when "10" & x"4b5" => DATA <= x"bebf";
            when "10" & x"4b6" => DATA <= x"c720";
            when "10" & x"4b7" => DATA <= x"0009";
            when "10" & x"4b8" => DATA <= x"4408";
            when "10" & x"4b9" => DATA <= x"ff33";
            when "10" & x"4ba" => DATA <= x"3ff8";
            when "10" & x"4bb" => DATA <= x"0124";
            when "10" & x"4bc" => DATA <= x"88ef";
            when "10" & x"4bd" => DATA <= x"f03d";
            when "10" & x"4be" => DATA <= x"0001";
            when "10" & x"4bf" => DATA <= x"03fd";
            when "10" & x"4c0" => DATA <= x"fe5e";
            when "10" & x"4c1" => DATA <= x"603f";
            when "10" & x"4c2" => DATA <= x"00ca";
            when "10" & x"4c3" => DATA <= x"07fb";
            when "10" & x"4c4" => DATA <= x"bdfe";
            when "10" & x"4c5" => DATA <= x"f079";
            when "10" & x"4c6" => DATA <= x"bfc1";
            when "10" & x"4c7" => DATA <= x"2f9e";
            when "10" & x"4c8" => DATA <= x"ff04";
            when "10" & x"4c9" => DATA <= x"805f";
            when "10" & x"4ca" => DATA <= x"e009";
            when "10" & x"4cb" => DATA <= x"ff00";
            when "10" & x"4cc" => DATA <= x"3f2f";
            when "10" & x"4cd" => DATA <= x"fc00";
            when "10" & x"4ce" => DATA <= x"0f7f";
            when "10" & x"4cf" => DATA <= x"a067";
            when "10" & x"4d0" => DATA <= x"fc00";
            when "10" & x"4d1" => DATA <= x"fc7f";
            when "10" & x"4d2" => DATA <= x"80e7";
            when "10" & x"4d3" => DATA <= x"fc01";
            when "10" & x"4d4" => DATA <= x"5fe0";
            when "10" & x"4d5" => DATA <= x"02a7";
            when "10" & x"4d6" => DATA <= x"7f80";
            when "10" & x"4d7" => DATA <= x"2bfc";
            when "10" & x"4d8" => DATA <= x"24ed";
            when "10" & x"4d9" => DATA <= x"eff7";
            when "10" & x"4da" => DATA <= x"01f9";
            when "10" & x"4db" => DATA <= x"fe00";
            when "10" & x"4dc" => DATA <= x"dff7";
            when "10" & x"4dd" => DATA <= x"e3fd";
            when "10" & x"4de" => DATA <= x"fdbf";
            when "10" & x"4df" => DATA <= x"ef17";
            when "10" & x"4e0" => DATA <= x"f807";
            when "10" & x"4e1" => DATA <= x"7fde";
            when "10" & x"4e2" => DATA <= x"eff0";
            when "10" & x"4e3" => DATA <= x"3cff";
            when "10" & x"4e4" => DATA <= x"a5df";
            when "10" & x"4e5" => DATA <= x"c4f2";
            when "10" & x"4e6" => DATA <= x"023f";
            when "10" & x"4e7" => DATA <= x"bfdd";
            when "10" & x"4e8" => DATA <= x"e000";
            when "10" & x"4e9" => DATA <= x"3281";
            when "10" & x"4ea" => DATA <= x"31df";
            when "10" & x"4eb" => DATA <= x"e087";
            when "10" & x"4ec" => DATA <= x"0200";
            when "10" & x"4ed" => DATA <= x"0a80";
            when "10" & x"4ee" => DATA <= x"eff4";
            when "10" & x"4ef" => DATA <= x"c3fd";
            when "10" & x"4f0" => DATA <= x"1e09";
            when "10" & x"4f1" => DATA <= x"20f7";
            when "10" & x"4f2" => DATA <= x"f801";
            when "10" & x"4f3" => DATA <= x"fe6d";
            when "10" & x"4f4" => DATA <= x"1220";
            when "10" & x"4f5" => DATA <= x"3bfc";
            when "10" & x"4f6" => DATA <= x"007f";
            when "10" & x"4f7" => DATA <= x"0005";
            when "10" & x"4f8" => DATA <= x"166d";
            when "10" & x"4f9" => DATA <= x"b7eb";
            when "10" & x"4fa" => DATA <= x"fc00";
            when "10" & x"4fb" => DATA <= x"f878";
            when "10" & x"4fc" => DATA <= x"1027";
            when "10" & x"4fd" => DATA <= x"fde0";
            when "10" & x"4fe" => DATA <= x"ff28";
            when "10" & x"4ff" => DATA <= x"9827";
            when "10" & x"500" => DATA <= x"fc38";
            when "10" & x"501" => DATA <= x"df77";
            when "10" & x"502" => DATA <= x"8413";
            when "10" & x"503" => DATA <= x"e6fa";
            when "10" & x"504" => DATA <= x"ff00";
            when "10" & x"505" => DATA <= x"d7fb";
            when "10" & x"506" => DATA <= x"ac01";
            when "10" & x"507" => DATA <= x"dfe0";
            when "10" & x"508" => DATA <= x"03fb";
            when "10" & x"509" => DATA <= x"fc42";
            when "10" & x"50a" => DATA <= x"f0ef";
            when "10" & x"50b" => DATA <= x"f005";
            when "10" & x"50c" => DATA <= x"7f80";
            when "10" & x"50d" => DATA <= x"67fc";
            when "10" & x"50e" => DATA <= x"000f";
            when "10" & x"50f" => DATA <= x"7780";
            when "10" & x"510" => DATA <= x"2b8c";
            when "10" & x"511" => DATA <= x"c6e3";
            when "10" & x"512" => DATA <= x"7628";
            when "10" & x"513" => DATA <= x"07e4";
            when "10" & x"514" => DATA <= x"0793";
            when "10" & x"515" => DATA <= x"e5e3";
            when "10" & x"516" => DATA <= x"5f8f";
            when "10" & x"517" => DATA <= x"f703";
            when "10" & x"518" => DATA <= x"fedf";
            when "10" & x"519" => DATA <= x"dfe7";
            when "10" & x"51a" => DATA <= x"f432";
            when "10" & x"51b" => DATA <= x"2aa7";
            when "10" & x"51c" => DATA <= x"9ed5";
            when "10" & x"51d" => DATA <= x"fe40";
            when "10" & x"51e" => DATA <= x"fff0";
            when "10" & x"51f" => DATA <= x"05ff";
            when "10" & x"520" => DATA <= x"bb40";
            when "10" & x"521" => DATA <= x"085e";
            when "10" & x"522" => DATA <= x"ff16";
            when "10" & x"523" => DATA <= x"229f";
            when "10" & x"524" => DATA <= x"e100";
            when "10" & x"525" => DATA <= x"e77f";
            when "10" & x"526" => DATA <= x"8007";
            when "10" & x"527" => DATA <= x"effa";
            when "10" & x"528" => DATA <= x"00ae";
            when "10" & x"529" => DATA <= x"f7f8";
            when "10" & x"52a" => DATA <= x"107c";
            when "10" & x"52b" => DATA <= x"ff00";
            when "10" & x"52c" => DATA <= x"27bb";
            when "10" & x"52d" => DATA <= x"fc00";
            when "10" & x"52e" => DATA <= x"e27f";
            when "10" & x"52f" => DATA <= x"800b";
            when "10" & x"530" => DATA <= x"9dfe";
            when "10" & x"531" => DATA <= x"c047";
            when "10" & x"532" => DATA <= x"bfe8";
            when "10" & x"533" => DATA <= x"01b6";
            when "10" & x"534" => DATA <= x"df7f";
            when "10" & x"535" => DATA <= x"8011";
            when "10" & x"536" => DATA <= x"eff0";
            when "10" & x"537" => DATA <= x"008b";
            when "10" & x"538" => DATA <= x"bfc2";
            when "10" & x"539" => DATA <= x"0e77";
            when "10" & x"53a" => DATA <= x"f801";
            when "10" & x"53b" => DATA <= x"80f7";
            when "10" & x"53c" => DATA <= x"aff0";
            when "10" & x"53d" => DATA <= x"057f";
            when "10" & x"53e" => DATA <= x"8027";
            when "10" & x"53f" => DATA <= x"fd78";
            when "10" & x"540" => DATA <= x"033f";
            when "10" & x"541" => DATA <= x"8800";
            when "10" & x"542" => DATA <= x"6efa";
            when "10" & x"543" => DATA <= x"ff0b";
            when "10" & x"544" => DATA <= x"8807";
            when "10" & x"545" => DATA <= x"8602";
            when "10" & x"546" => DATA <= x"377f";
            when "10" & x"547" => DATA <= x"9e5e";
            when "10" & x"548" => DATA <= x"2491";
            when "10" & x"549" => DATA <= x"405f";
            when "10" & x"54a" => DATA <= x"bfc8";
            when "10" & x"54b" => DATA <= x"0df0";
            when "10" & x"54c" => DATA <= x"d180";
            when "10" & x"54d" => DATA <= x"80fb";
            when "10" & x"54e" => DATA <= x"7bbf";
            when "10" & x"54f" => DATA <= x"c700";
            when "10" & x"550" => DATA <= x"05b8";
            when "10" & x"551" => DATA <= x"f810";
            when "10" & x"552" => DATA <= x"ff7b";
            when "10" & x"553" => DATA <= x"bfeb";
            when "10" & x"554" => DATA <= x"f1fa";
            when "10" & x"555" => DATA <= x"f104";
            when "10" & x"556" => DATA <= x"3eeb";
            when "10" & x"557" => DATA <= x"fc86";
            when "10" & x"558" => DATA <= x"e30b";
            when "10" & x"559" => DATA <= x"88c6";
            when "10" & x"55a" => DATA <= x"03fa";
            when "10" & x"55b" => DATA <= x"ff40";
            when "10" & x"55c" => DATA <= x"2051";
            when "10" & x"55d" => DATA <= x"0002";
            when "10" & x"55e" => DATA <= x"0143";
            when "10" & x"55f" => DATA <= x"5381";
            when "10" & x"560" => DATA <= x"ddb9";
            when "10" & x"561" => DATA <= x"bbff";
            when "10" & x"562" => DATA <= x"eef7";
            when "10" & x"563" => DATA <= x"f713";
            when "10" & x"564" => DATA <= x"8f0e";
            when "10" & x"565" => DATA <= x"0783";
            when "10" & x"566" => DATA <= x"81e0";
            when "10" & x"567" => DATA <= x"e07b";
            when "10" & x"568" => DATA <= x"bff7";
            when "10" & x"569" => DATA <= x"bd1e";
            when "10" & x"56a" => DATA <= x"ef7f";
            when "10" & x"56b" => DATA <= x"87a7";
            when "10" & x"56c" => DATA <= x"f802";
            when "10" & x"56d" => DATA <= x"3f7f";
            when "10" & x"56e" => DATA <= x"d000";
            when "10" & x"56f" => DATA <= x"042a";
            when "10" & x"570" => DATA <= x"0138";
            when "10" & x"571" => DATA <= x"0001";
            when "10" & x"572" => DATA <= x"fc00";
            when "10" & x"573" => DATA <= x"1000";
            when "10" & x"574" => DATA <= x"382b";
            when "10" & x"575" => DATA <= x"c2b8";
            when "10" & x"576" => DATA <= x"11ca";
            when "10" & x"577" => DATA <= x"8570";
            when "10" & x"578" => DATA <= x"fcff";
            when "10" & x"579" => DATA <= x"47ef";
            when "10" & x"57a" => DATA <= x"f3fb";
            when "10" & x"57b" => DATA <= x"fdbe";
            when "10" & x"57c" => DATA <= x"0106";
            when "10" & x"57d" => DATA <= x"b841";
            when "10" & x"57e" => DATA <= x"2e13";
            when "10" & x"57f" => DATA <= x"d9f0";
            when "10" & x"580" => DATA <= x"e080";
            when "10" & x"581" => DATA <= x"000f";
            when "10" & x"582" => DATA <= x"d00c";
            when "10" & x"583" => DATA <= x"f07d";
            when "10" & x"584" => DATA <= x"0e81";
            when "10" & x"585" => DATA <= x"0004";
            when "10" & x"586" => DATA <= x"976b";
            when "10" & x"587" => DATA <= x"ff80";
            when "10" & x"588" => DATA <= x"0400";
            when "10" & x"589" => DATA <= x"04d2";
            when "10" & x"58a" => DATA <= x"7dbe";
            when "10" & x"58b" => DATA <= x"c040";
            when "10" & x"58c" => DATA <= x"0018";
            when "10" & x"58d" => DATA <= x"a216";
            when "10" & x"58e" => DATA <= x"8079";
            when "10" & x"58f" => DATA <= x"eefd";
            when "10" & x"590" => DATA <= x"003f";
            when "10" & x"591" => DATA <= x"4400";
            when "10" & x"592" => DATA <= x"1028";
            when "10" & x"593" => DATA <= x"02bf";
            when "10" & x"594" => DATA <= x"dc0f";
            when "10" & x"595" => DATA <= x"f102";
            when "10" & x"596" => DATA <= x"49e0";
            when "10" & x"597" => DATA <= x"007f";
            when "10" & x"598" => DATA <= x"bdc0";
            when "10" & x"599" => DATA <= x"6ff0";
            when "10" & x"59a" => DATA <= x"0010";
            when "10" & x"59b" => DATA <= x"3e80";
            when "10" & x"59c" => DATA <= x"6f87";
            when "10" & x"59d" => DATA <= x"d80b";
            when "10" & x"59e" => DATA <= x"f400";
            when "10" & x"59f" => DATA <= x"0800";
            when "10" & x"5a0" => DATA <= x"8069";
            when "10" & x"5a1" => DATA <= x"91c0";
            when "10" & x"5a2" => DATA <= x"2fc0";
            when "10" & x"5a3" => DATA <= x"2000";
            when "10" & x"5a4" => DATA <= x"915f";
            when "10" & x"5a5" => DATA <= x"e125";
            when "10" & x"5a6" => DATA <= x"2010";
            when "10" & x"5a7" => DATA <= x"4140";
            when "10" & x"5a8" => DATA <= x"15fe";
            when "10" & x"5a9" => DATA <= x"0912";
            when "10" & x"5aa" => DATA <= x"8808";
            when "10" & x"5ab" => DATA <= x"a047";
            when "10" & x"5ac" => DATA <= x"e08d";
            when "10" & x"5ad" => DATA <= x"86fe";
            when "10" & x"5ae" => DATA <= x"023c";
            when "10" & x"5af" => DATA <= x"0442";
            when "10" & x"5b0" => DATA <= x"10f8";
            when "10" & x"5b1" => DATA <= x"02bf";
            when "10" & x"5b2" => DATA <= x"d80f";
            when "10" & x"5b3" => DATA <= x"f422";
            when "10" & x"5b4" => DATA <= x"01dc";
            when "10" & x"5b5" => DATA <= x"0171";
            when "10" & x"5b6" => DATA <= x"bbc1";
            when "10" & x"5b7" => DATA <= x"eff0";
            when "10" & x"5b8" => DATA <= x"8090";
            when "10" & x"5b9" => DATA <= x"fe00";
            when "10" & x"5ba" => DATA <= x"5f9f";
            when "10" & x"5bb" => DATA <= x"d007";
            when "10" & x"5bc" => DATA <= x"fa00";
            when "10" & x"5bd" => DATA <= x"42ba";
            when "10" & x"5be" => DATA <= x"80cc";
            when "10" & x"5bf" => DATA <= x"6038";
            when "10" & x"5c0" => DATA <= x"f091";
            when "10" & x"5c1" => DATA <= x"400f";
            when "10" & x"5c2" => DATA <= x"f003";
            when "10" & x"5c3" => DATA <= x"fc96";
            when "10" & x"5c4" => DATA <= x"48a0";
            when "10" & x"5c5" => DATA <= x"0121";
            when "10" & x"5c6" => DATA <= x"fd80";
            when "10" & x"5c7" => DATA <= x"9f09";
            when "10" & x"5c8" => DATA <= x"0005";
            when "10" & x"5c9" => DATA <= x"4ca7";
            when "10" & x"5ca" => DATA <= x"f061";
            when "10" & x"5cb" => DATA <= x"e2ff";
            when "10" & x"5cc" => DATA <= x"013f";
            when "10" & x"5cd" => DATA <= x"0a25";
            when "10" & x"5ce" => DATA <= x"023a";
            when "10" & x"5cf" => DATA <= x"12bf";
            when "10" & x"5d0" => DATA <= x"dc0f";
            when "10" & x"5d1" => DATA <= x"f311";
            when "10" & x"5d2" => DATA <= x"01fc";
            when "10" & x"5d3" => DATA <= x"0079";
            when "10" & x"5d4" => DATA <= x"3ec1";
            when "10" & x"5d5" => DATA <= x"6ff0";
            when "10" & x"5d6" => DATA <= x"5825";
            when "10" & x"5d7" => DATA <= x"be80";
            when "10" & x"5d8" => DATA <= x"0f97";
            when "10" & x"5d9" => DATA <= x"c801";
            when "10" & x"5da" => DATA <= x"fa00";
            when "10" & x"5db" => DATA <= x"01bc";
            when "10" & x"5dc" => DATA <= x"002f";
            when "10" & x"5dd" => DATA <= x"1008";
            when "10" & x"5de" => DATA <= x"fc10";
            when "10" & x"5df" => DATA <= x"0040";
            when "10" & x"5e0" => DATA <= x"3fc0";
            when "10" & x"5e1" => DATA <= x"0ffa";
            when "10" & x"5e2" => DATA <= x"4900";
            when "10" & x"5e3" => DATA <= x"2004";
            when "10" & x"5e4" => DATA <= x"80f4";
            when "10" & x"5e5" => DATA <= x"02dd";
            when "10" & x"5e6" => DATA <= x"06c0";
            when "10" & x"5e7" => DATA <= x"0404";
            when "10" & x"5e8" => DATA <= x"0483";
            when "10" & x"5e9" => DATA <= x"a003";
            when "10" & x"5ea" => DATA <= x"fc00";
            when "10" & x"5eb" => DATA <= x"ffa0";
            when "10" & x"5ec" => DATA <= x"4003";
            when "10" & x"5ed" => DATA <= x"f400";
            when "10" & x"5ee" => DATA <= x"ff40";
            when "10" & x"5ef" => DATA <= x"bfc0";
            when "10" & x"5f0" => DATA <= x"66c3";
            when "10" & x"5f1" => DATA <= x"4bfc";
            when "10" & x"5f2" => DATA <= x"00ff";
            when "10" & x"5f3" => DATA <= x"04bf";
            when "10" & x"5f4" => DATA <= x"c014";
            when "10" & x"5f5" => DATA <= x"02ff";
            when "10" & x"5f6" => DATA <= x"0036";
            when "10" & x"5f7" => DATA <= x"c386";
            when "10" & x"5f8" => DATA <= x"3085";
            when "10" & x"5f9" => DATA <= x"003f";
            when "10" & x"5fa" => DATA <= x"c00f";
            when "10" & x"5fb" => DATA <= x"f480";
            when "10" & x"5fc" => DATA <= x"4840";
            when "10" & x"5fd" => DATA <= x"0024";
            when "10" & x"5fe" => DATA <= x"87c0";
            when "10" & x"5ff" => DATA <= x"0770";
            when "10" & x"600" => DATA <= x"3201";
            when "10" & x"601" => DATA <= x"6021";
            when "10" & x"602" => DATA <= x"241d";
            when "10" & x"603" => DATA <= x"002f";
            when "10" & x"604" => DATA <= x"f00b";
            when "10" & x"605" => DATA <= x"fc10";
            when "10" & x"606" => DATA <= x"2830";
            when "10" & x"607" => DATA <= x"3e80";
            when "10" & x"608" => DATA <= x"0ff0";
            when "10" & x"609" => DATA <= x"03fc";
            when "10" & x"60a" => DATA <= x"0d5b";
            when "10" & x"60b" => DATA <= x"0ff0";
            when "10" & x"60c" => DATA <= x"03fc";
            when "10" & x"60d" => DATA <= x"20ff";
            when "10" & x"60e" => DATA <= x"2050";
            when "10" & x"60f" => DATA <= x"13fd";
            when "10" & x"610" => DATA <= x"e037";
            when "10" & x"611" => DATA <= x"7031";
            when "10" & x"612" => DATA <= x"c802";
            when "10" & x"613" => DATA <= x"0401";
            when "10" & x"614" => DATA <= x"4dfe";
            when "10" & x"615" => DATA <= x"fd7f";
            when "10" & x"616" => DATA <= x"00d0";
            when "10" & x"617" => DATA <= x"04b0";
            when "10" & x"618" => DATA <= x"0015";
            when "10" & x"619" => DATA <= x"fc3e";
            when "10" & x"61a" => DATA <= x"7f80";
            when "10" & x"61b" => DATA <= x"1108";
            when "10" & x"61c" => DATA <= x"200b";
            when "10" & x"61d" => DATA <= x"c0fe";
            when "10" & x"61e" => DATA <= x"fd7f";
            when "10" & x"61f" => DATA <= x"d000";
            when "10" & x"620" => DATA <= x"4804";
            when "10" & x"621" => DATA <= x"bfa7";
            when "10" & x"622" => DATA <= x"e7fd";
            when "10" & x"623" => DATA <= x"000c";
            when "10" & x"624" => DATA <= x"8104";
            when "10" & x"625" => DATA <= x"2eff";
            when "10" & x"626" => DATA <= x"0010";
            when "10" & x"627" => DATA <= x"08a0";
            when "10" & x"628" => DATA <= x"0600";
            when "10" & x"629" => DATA <= x"1ebf";
            when "10" & x"62a" => DATA <= x"c006";
            when "10" & x"62b" => DATA <= x"c6a2";
            when "10" & x"62c" => DATA <= x"113c";
            when "10" & x"62d" => DATA <= x"8e5f";
            when "10" & x"62e" => DATA <= x"bfc0";
            when "10" & x"62f" => DATA <= x"15fd";
            when "10" & x"630" => DATA <= x"dfef";
            when "10" & x"631" => DATA <= x"77f8";
            when "10" & x"632" => DATA <= x"02bf";
            when "10" & x"633" => DATA <= x"e401";
            when "10" & x"634" => DATA <= x"f000";
            when "10" & x"635" => DATA <= x"aff0";
            when "10" & x"636" => DATA <= x"03f1";
            when "10" & x"637" => DATA <= x"181c";
            when "10" & x"638" => DATA <= x"3e9f";
            when "10" & x"639" => DATA <= x"2bfd";
            when "10" & x"63a" => DATA <= x"e1de";
            when "10" & x"63b" => DATA <= x"35e6";
            when "10" & x"63c" => DATA <= x"ef9f";
            when "10" & x"63d" => DATA <= x"f638";
            when "10" & x"63e" => DATA <= x"1d4f";
            when "10" & x"63f" => DATA <= x"3fef";
            when "10" & x"640" => DATA <= x"47b0";
            when "10" & x"641" => DATA <= x"01e6";
            when "10" & x"642" => DATA <= x"f7ef";
            when "10" & x"643" => DATA <= x"f773";
            when "10" & x"644" => DATA <= x"fc00";
            when "10" & x"645" => DATA <= x"2e97";
            when "10" & x"646" => DATA <= x"f3d8";
            when "10" & x"647" => DATA <= x"8068";
            when "10" & x"648" => DATA <= x"3e6c";
            when "10" & x"649" => DATA <= x"a048";
            when "10" & x"64a" => DATA <= x"a016";
            when "10" & x"64b" => DATA <= x"2916";
            when "10" & x"64c" => DATA <= x"8159";
            when "10" & x"64d" => DATA <= x"4404";
            when "10" & x"64e" => DATA <= x"1761";
            when "10" & x"64f" => DATA <= x"d001";
            when "10" & x"650" => DATA <= x"cc00";
            when "10" & x"651" => DATA <= x"2011";
            when "10" & x"652" => DATA <= x"0c82";
            when "10" & x"653" => DATA <= x"4800";
            when "10" & x"654" => DATA <= x"011c";
            when "10" & x"655" => DATA <= x"8642";
            when "10" & x"656" => DATA <= x"1988";
            when "10" & x"657" => DATA <= x"d064";
            when "10" & x"658" => DATA <= x"33fa";
            when "10" & x"659" => DATA <= x"fdd0";
            when "10" & x"65a" => DATA <= x"0401";
            when "10" & x"65b" => DATA <= x"5000";
            when "10" & x"65c" => DATA <= x"a000";
            when "10" & x"65d" => DATA <= x"ff09";
            when "10" & x"65e" => DATA <= x"8001";
            when "10" & x"65f" => DATA <= x"286e";
            when "10" & x"660" => DATA <= x"003f";
            when "10" & x"661" => DATA <= x"8424";
            when "10" & x"662" => DATA <= x"0100";
            when "10" & x"663" => DATA <= x"005f";
            when "10" & x"664" => DATA <= x"0040";
            when "10" & x"665" => DATA <= x"802a";
            when "10" & x"666" => DATA <= x"0009";
            when "10" & x"667" => DATA <= x"8315";
            when "10" & x"668" => DATA <= x"ebc0";
            when "10" & x"669" => DATA <= x"0200";
            when "10" & x"66a" => DATA <= x"0208";
            when "10" & x"66b" => DATA <= x"1002";
            when "10" & x"66c" => DATA <= x"1c41";
            when "10" & x"66d" => DATA <= x"5100";
            when "10" & x"66e" => DATA <= x"0400";
            when "10" & x"66f" => DATA <= x"0ca4";
            when "10" & x"670" => DATA <= x"07cb";
            when "10" & x"671" => DATA <= x"3240";
            when "10" & x"672" => DATA <= x"0440";
            when "10" & x"673" => DATA <= x"12c1";
            when "10" & x"674" => DATA <= x"e840";
            when "10" & x"675" => DATA <= x"0fa8";
            when "10" & x"676" => DATA <= x"0000";
            when "10" & x"677" => DATA <= x"81b6";
            when "10" & x"678" => DATA <= x"9068";
            when "10" & x"679" => DATA <= x"07d8";
            when "10" & x"67a" => DATA <= x"1480";
            when "10" & x"67b" => DATA <= x"c0a0";
            when "10" & x"67c" => DATA <= x"0418";
            when "10" & x"67d" => DATA <= x"000e";
            when "10" & x"67e" => DATA <= x"a069";
            when "10" & x"67f" => DATA <= x"01dc";
            when "10" & x"680" => DATA <= x"0617";
            when "10" & x"681" => DATA <= x"1380";
            when "10" & x"682" => DATA <= x"c062";
            when "10" & x"683" => DATA <= x"0138";
            when "10" & x"684" => DATA <= x"2801";
            when "10" & x"685" => DATA <= x"00f0";
            when "10" & x"686" => DATA <= x"002c";
            when "10" & x"687" => DATA <= x"57cf";
            when "10" & x"688" => DATA <= x"4afc";
            when "10" & x"689" => DATA <= x"7a3e";
            when "10" & x"68a" => DATA <= x"5f8f";
            when "10" & x"68b" => DATA <= x"d7cb";
            when "10" & x"68c" => DATA <= x"d026";
            when "10" & x"68d" => DATA <= x"0311";
            when "10" & x"68e" => DATA <= x"81e8";
            when "10" & x"68f" => DATA <= x"5e81";
            when "10" & x"690" => DATA <= x"d88c";
            when "10" & x"691" => DATA <= x"0702";
            when "10" & x"692" => DATA <= x"0120";
            when "10" & x"693" => DATA <= x"d000";
            when "10" & x"694" => DATA <= x"0101";
            when "10" & x"695" => DATA <= x"c0da";
            when "10" & x"696" => DATA <= x"0c7f";
            when "10" & x"697" => DATA <= x"3e2b";
            when "10" & x"698" => DATA <= x"f9bf";
            when "10" & x"699" => DATA <= x"5ffb";
            when "10" & x"69a" => DATA <= x"bef7";
            when "10" & x"69b" => DATA <= x"affd";
            when "10" & x"69c" => DATA <= x"f718";
            when "10" & x"69d" => DATA <= x"db88";
            when "10" & x"69e" => DATA <= x"0687";
            when "10" & x"69f" => DATA <= x"a870";
            when "10" & x"6a0" => DATA <= x"3d43";
            when "10" & x"6a1" => DATA <= x"81ee";
            when "10" & x"6a2" => DATA <= x"efaf";
            when "10" & x"6a3" => DATA <= x"feef";
            when "10" & x"6a4" => DATA <= x"afe7";
            when "10" & x"6a5" => DATA <= x"b3dd";
            when "10" & x"6a6" => DATA <= x"ff5f";
            when "10" & x"6a7" => DATA <= x"c7e0";
            when "10" & x"6a8" => DATA <= x"0944";
            when "10" & x"6a9" => DATA <= x"2271";
            when "10" & x"6aa" => DATA <= x"0880";
            when "10" & x"6ab" => DATA <= x"4a74";
            when "10" & x"6ac" => DATA <= x"0010";
            when "10" & x"6ad" => DATA <= x"0008";
            when "10" & x"6ae" => DATA <= x"000f";
            when "10" & x"6af" => DATA <= x"c408";
            when "10" & x"6b0" => DATA <= x"0114";
            when "10" & x"6b1" => DATA <= x"8202";
            when "10" & x"6b2" => DATA <= x"5043";
            when "10" & x"6b3" => DATA <= x"0102";
            when "10" & x"6b4" => DATA <= x"807e";
            when "10" & x"6b5" => DATA <= x"aff7";
            when "10" & x"6b6" => DATA <= x"fdfa";
            when "10" & x"6b7" => DATA <= x"7c3c";
            when "10" & x"6b8" => DATA <= x"804c";
            when "10" & x"6b9" => DATA <= x"3cf8";
            when "10" & x"6ba" => DATA <= x"fc4e";
            when "10" & x"6bb" => DATA <= x"87c3";
            when "10" & x"6bc" => DATA <= x"c5d4";
            when "10" & x"6bd" => DATA <= x"e8f4";
            when "10" & x"6be" => DATA <= x"3a4d";
            when "10" & x"6bf" => DATA <= x"0250";
            when "10" & x"6c0" => DATA <= x"0121";
            when "10" & x"6c1" => DATA <= x"fef4";
            when "10" & x"6c2" => DATA <= x"1300";
            when "10" & x"6c3" => DATA <= x"b801";
            when "10" & x"6c4" => DATA <= x"04ff";
            when "10" & x"6c5" => DATA <= x"0200";
            when "10" & x"6c6" => DATA <= x"01ef";
            when "10" & x"6c7" => DATA <= x"c7e8";
            when "10" & x"6c8" => DATA <= x"0400";
            when "10" & x"6c9" => DATA <= x"eb00";
            when "10" & x"6ca" => DATA <= x"200f";
            when "10" & x"6cb" => DATA <= x"55ff";
            when "10" & x"6cc" => DATA <= x"400f";
            when "10" & x"6cd" => DATA <= x"f3a0";
            when "10" & x"6ce" => DATA <= x"e4d1";
            when "10" & x"6cf" => DATA <= x"5fe0";
            when "10" & x"6d0" => DATA <= x"1003";
            when "10" & x"6d1" => DATA <= x"fc02";
            when "10" & x"6d2" => DATA <= x"3101";
            when "10" & x"6d3" => DATA <= x"07d7";
            when "10" & x"6d4" => DATA <= x"e800";
            when "10" & x"6d5" => DATA <= x"03fd";
            when "10" & x"6d6" => DATA <= x"34da";
            when "10" & x"6d7" => DATA <= x"003f";
            when "10" & x"6d8" => DATA <= x"29f0";
            when "10" & x"6d9" => DATA <= x"faff";
            when "10" & x"6da" => DATA <= x"a010";
            when "10" & x"6db" => DATA <= x"8013";
            when "10" & x"6dc" => DATA <= x"801f";
            when "10" & x"6dd" => DATA <= x"f400";
            when "10" & x"6de" => DATA <= x"2a90";
            when "10" & x"6df" => DATA <= x"07fd";
            when "10" & x"6e0" => DATA <= x"002c";
            when "10" & x"6e1" => DATA <= x"9f55";
            when "10" & x"6e2" => DATA <= x"f0a0";
            when "10" & x"6e3" => DATA <= x"7f80";
            when "10" & x"6e4" => DATA <= x"0085";
            when "10" & x"6e5" => DATA <= x"3eff";
            when "10" & x"6e6" => DATA <= x"3f3f";
            when "10" & x"6e7" => DATA <= x"c002";
            when "10" & x"6e8" => DATA <= x"627e";
            when "10" & x"6e9" => DATA <= x"ffd1";
            when "10" & x"6ea" => DATA <= x"c0bf";
            when "10" & x"6eb" => DATA <= x"9fcd";
            when "10" & x"6ec" => DATA <= x"aff0";
            when "10" & x"6ed" => DATA <= x"0004";
            when "10" & x"6ee" => DATA <= x"0039";
            when "10" & x"6ef" => DATA <= x"1c2e";
            when "10" & x"6f0" => DATA <= x"178e";
            when "10" & x"6f1" => DATA <= x"f7f1";
            when "10" & x"6f2" => DATA <= x"f800";
            when "10" & x"6f3" => DATA <= x"08e0";
            when "10" & x"6f4" => DATA <= x"07fb";
            when "10" & x"6f5" => DATA <= x"e400";
            when "10" & x"6f6" => DATA <= x"7090";
            when "10" & x"6f7" => DATA <= x"07f8";
            when "10" & x"6f8" => DATA <= x"0008";
            when "10" & x"6f9" => DATA <= x"067e";
            when "10" & x"6fa" => DATA <= x"d7e2";
            when "10" & x"6fb" => DATA <= x"a9f2";
            when "10" & x"6fc" => DATA <= x"ff07";
            when "10" & x"6fd" => DATA <= x"803b";
            when "10" & x"6fe" => DATA <= x"fd54";
            when "10" & x"6ff" => DATA <= x"d77f";
            when "10" & x"700" => DATA <= x"d007";
            when "10" & x"701" => DATA <= x"7faa";
            when "10" & x"702" => DATA <= x"abfe";
            when "10" & x"703" => DATA <= x"8017";
            when "10" & x"704" => DATA <= x"f47e";
            when "10" & x"705" => DATA <= x"2aaf";
            when "10" & x"706" => DATA <= x"fa00";
            when "10" & x"707" => DATA <= x"e3c6";
            when "10" & x"708" => DATA <= x"e870";
            when "10" & x"709" => DATA <= x"3fa0";
            when "10" & x"70a" => DATA <= x"0ffa";
            when "10" & x"70b" => DATA <= x"80a0";
            when "10" & x"70c" => DATA <= x"0403";
            when "10" & x"70d" => DATA <= x"0010";
            when "10" & x"70e" => DATA <= x"ff00";
            when "10" & x"70f" => DATA <= x"0fc0";
            when "10" & x"710" => DATA <= x"0c07";
            when "10" & x"711" => DATA <= x"fafc";
            when "10" & x"712" => DATA <= x"00ff";
            when "10" & x"713" => DATA <= x"003f";
            when "10" & x"714" => DATA <= x"0c15";
            when "10" & x"715" => DATA <= x"fefb";
            when "10" & x"716" => DATA <= x"003f";
            when "10" & x"717" => DATA <= x"c00f";
            when "10" & x"718" => DATA <= x"f77f";
            when "10" & x"719" => DATA <= x"7f80";
            when "10" & x"71a" => DATA <= x"1fe0";
            when "10" & x"71b" => DATA <= x"0eff";
            when "10" & x"71c" => DATA <= x"2590";
            when "10" & x"71d" => DATA <= x"ca0f";
            when "10" & x"71e" => DATA <= x"f003";
            when "10" & x"71f" => DATA <= x"fdbe";
            when "10" & x"720" => DATA <= x"ffe0";
            when "10" & x"721" => DATA <= x"07f8";
            when "10" & x"722" => DATA <= x"01fe";
            when "10" & x"723" => DATA <= x"f37f";
            when "10" & x"724" => DATA <= x"8828";
            when "10" & x"725" => DATA <= x"01fe";
            when "10" & x"726" => DATA <= x"007f";
            when "10" & x"727" => DATA <= x"8045";
            when "10" & x"728" => DATA <= x"35fe";
            when "10" & x"729" => DATA <= x"007f";
            when "10" & x"72a" => DATA <= x"801f";
            when "10" & x"72b" => DATA <= x"e115";
            when "10" & x"72c" => DATA <= x"abfc";
            when "10" & x"72d" => DATA <= x"fe00";
            when "10" & x"72e" => DATA <= x"7f80";
            when "10" & x"72f" => DATA <= x"1fe0";
            when "10" & x"730" => DATA <= x"04f5";
            when "10" & x"731" => DATA <= x"7f80";
            when "10" & x"732" => DATA <= x"1fe0";
            when "10" & x"733" => DATA <= x"0038";
            when "10" & x"734" => DATA <= x"01fc";
            when "10" & x"735" => DATA <= x"1343";
            when "10" & x"736" => DATA <= x"a81f";
            when "10" & x"737" => DATA <= x"f400";
            when "10" & x"738" => DATA <= x"c67f";
            when "10" & x"739" => DATA <= x"82e8";
            when "10" & x"73a" => DATA <= x"0c46";
            when "10" & x"73b" => DATA <= x"1800";
            when "10" & x"73c" => DATA <= x"0e47";
            when "10" & x"73d" => DATA <= x"e005";
            when "10" & x"73e" => DATA <= x"00e2";
            when "10" & x"73f" => DATA <= x"8004";
            when "10" & x"740" => DATA <= x"0030";
            when "10" & x"741" => DATA <= x"1001";
            when "10" & x"742" => DATA <= x"d4ff";
            when "10" & x"743" => DATA <= x"a001";
            when "10" & x"744" => DATA <= x"1700";
            when "10" & x"745" => DATA <= x"17cf";
            when "10" & x"746" => DATA <= x"e002";
            when "10" & x"747" => DATA <= x"028b";
            when "10" & x"748" => DATA <= x"8000";
            when "10" & x"749" => DATA <= x"6e00";
            when "10" & x"74a" => DATA <= x"a0d0";
            when "10" & x"74b" => DATA <= x"409e";
            when "10" & x"74c" => DATA <= x"2180";
            when "10" & x"74d" => DATA <= x"0f6b";
            when "10" & x"74e" => DATA <= x"9582";
            when "10" & x"74f" => DATA <= x"ec30";
            when "10" & x"750" => DATA <= x"e750";
            when "10" & x"751" => DATA <= x"8017";
            when "10" & x"752" => DATA <= x"8fea";
            when "10" & x"753" => DATA <= x"fc1f";
            when "10" & x"754" => DATA <= x"2fdf";
            when "10" & x"755" => DATA <= x"e006";
            when "10" & x"756" => DATA <= x"bbfc";
            when "10" & x"757" => DATA <= x"4aff";
            when "10" & x"758" => DATA <= x"101e";
            when "10" & x"759" => DATA <= x"1fe0";
            when "10" & x"75a" => DATA <= x"069b";
            when "10" & x"75b" => DATA <= x"fc80";
            when "10" & x"75c" => DATA <= x"ff00";
            when "10" & x"75d" => DATA <= x"0d1f";
            when "10" & x"75e" => DATA <= x"e000";
            when "10" & x"75f" => DATA <= x"3bfc";
            when "10" & x"760" => DATA <= x"02ff";
            when "10" & x"761" => DATA <= x"0002";
            when "10" & x"762" => DATA <= x"07ef";
            when "10" & x"763" => DATA <= x"0af3";
            when "10" & x"764" => DATA <= x"793c";
            when "10" & x"765" => DATA <= x"de0f";
            when "10" & x"766" => DATA <= x"f415";
            when "10" & x"767" => DATA <= x"03d4";
            when "10" & x"768" => DATA <= x"381d";
            when "10" & x"769" => DATA <= x"0e3f";
            when "10" & x"76a" => DATA <= x"7f80";
            when "10" & x"76b" => DATA <= x"0580";
            when "10" & x"76c" => DATA <= x"e900";
            when "10" & x"76d" => DATA <= x"4080";
            when "10" & x"76e" => DATA <= x"0a25";
            when "10" & x"76f" => DATA <= x"0e00";
            when "10" & x"770" => DATA <= x"57be";
            when "10" & x"771" => DATA <= x"c00f";
            when "10" & x"772" => DATA <= x"65a0";
            when "10" & x"773" => DATA <= x"3280";
            when "10" & x"774" => DATA <= x"1e4f";
            when "10" & x"775" => DATA <= x"a02b";
            when "10" & x"776" => DATA <= x"8abf";
            when "10" & x"777" => DATA <= x"df00";
            when "10" & x"778" => DATA <= x"0038";
            when "10" & x"779" => DATA <= x"7c00";
            when "10" & x"77a" => DATA <= x"f7af";
            when "10" & x"77b" => DATA <= x"f378";
            when "10" & x"77c" => DATA <= x"01fe";
            when "10" & x"77d" => DATA <= x"8700";
            when "10" & x"77e" => DATA <= x"06ab";
            when "10" & x"77f" => DATA <= x"fc06";
            when "10" & x"780" => DATA <= x"f87f";
            when "10" & x"781" => DATA <= x"820e";
            when "10" & x"782" => DATA <= x"0749";
            when "10" & x"783" => DATA <= x"703f";
            when "10" & x"784" => DATA <= x"83d0";
            when "10" & x"785" => DATA <= x"e100";
            when "10" & x"786" => DATA <= x"03e0";
            when "10" & x"787" => DATA <= x"40bc";
            when "10" & x"788" => DATA <= x"5f00";
            when "10" & x"789" => DATA <= x"0600";
            when "10" & x"78a" => DATA <= x"0011";
            when "10" & x"78b" => DATA <= x"fca4";
            when "10" & x"78c" => DATA <= x"030a";
            when "10" & x"78d" => DATA <= x"5000";
            when "10" & x"78e" => DATA <= x"6800";
            when "10" & x"78f" => DATA <= x"1026";
            when "10" & x"790" => DATA <= x"0381";
            when "10" & x"791" => DATA <= x"f200";
            when "10" & x"792" => DATA <= x"8100";
            when "10" & x"793" => DATA <= x"2006";
            when "10" & x"794" => DATA <= x"eb92";
            when "10" & x"795" => DATA <= x"0500";
            when "10" & x"796" => DATA <= x"3c10";
            when "10" & x"797" => DATA <= x"0241";
            when "10" & x"798" => DATA <= x"100c";
            when "10" & x"799" => DATA <= x"0006";
            when "10" & x"79a" => DATA <= x"00d0";
            when "10" & x"79b" => DATA <= x"002c";
            when "10" & x"79c" => DATA <= x"4608";
            when "10" & x"79d" => DATA <= x"0094";
            when "10" & x"79e" => DATA <= x"4420";
            when "10" & x"79f" => DATA <= x"7389";
            when "10" & x"7a0" => DATA <= x"44e2";
            when "10" & x"7a1" => DATA <= x"f140";
            when "10" & x"7a2" => DATA <= x"0004";
            when "10" & x"7a3" => DATA <= x"8103";
            when "10" & x"7a4" => DATA <= x"8809";
            when "10" & x"7a5" => DATA <= x"1048";
            when "10" & x"7a6" => DATA <= x"0011";
            when "10" & x"7a7" => DATA <= x"9204";
            when "10" & x"7a8" => DATA <= x"e200";
            when "10" & x"7a9" => DATA <= x"001e";
            when "10" & x"7aa" => DATA <= x"4000";
            when "10" & x"7ab" => DATA <= x"30c0";
            when "10" & x"7ac" => DATA <= x"5400";
            when "10" & x"7ad" => DATA <= x"08a8";
            when "10" & x"7ae" => DATA <= x"2302";
            when "10" & x"7af" => DATA <= x"48c0";
            when "10" & x"7b0" => DATA <= x"9068";
            when "10" & x"7b1" => DATA <= x"001c";
            when "10" & x"7b2" => DATA <= x"0600";
            when "10" & x"7b3" => DATA <= x"0089";
            when "10" & x"7b4" => DATA <= x"c061";
            when "10" & x"7b5" => DATA <= x"5e28";
            when "10" & x"7b6" => DATA <= x"9f8f";
            when "10" & x"7b7" => DATA <= x"37e3";
            when "10" & x"7b8" => DATA <= x"c5e8";
            when "10" & x"7b9" => DATA <= x"7daf";
            when "10" & x"7ba" => DATA <= x"8743";
            when "10" & x"7bb" => DATA <= x"e02e";
            when "10" & x"7bc" => DATA <= x"d775";
            when "10" & x"7bd" => DATA <= x"a080";
            when "10" & x"7be" => DATA <= x"607a";
            when "10" & x"7bf" => DATA <= x"c752";
            when "10" & x"7c0" => DATA <= x"385e";
            when "10" & x"7c1" => DATA <= x"f400";
            when "10" & x"7c2" => DATA <= x"fe7f";
            when "10" & x"7c3" => DATA <= x"83df";
            when "10" & x"7c4" => DATA <= x"ce77";
            when "10" & x"7c5" => DATA <= x"fd00";
            when "10" & x"7c6" => DATA <= x"0040";
            when "10" & x"7c7" => DATA <= x"680e";
            when "10" & x"7c8" => DATA <= x"df2f";
            when "10" & x"7c9" => DATA <= x"80c0";
            when "10" & x"7ca" => DATA <= x"0d06";
            when "10" & x"7cb" => DATA <= x"fd7b";
            when "10" & x"7cc" => DATA <= x"81e8";
            when "10" & x"7cd" => DATA <= x"01f9";
            when "10" & x"7ce" => DATA <= x"5ee0";
            when "10" & x"7cf" => DATA <= x"1e00";
            when "10" & x"7d0" => DATA <= x"2073";
            when "10" & x"7d1" => DATA <= x"8d0e";
            when "10" & x"7d2" => DATA <= x"70f0";
            when "10" & x"7d3" => DATA <= x"7287";
            when "10" & x"7d4" => DATA <= x"afbe";
            when "10" & x"7d5" => DATA <= x"bfe7";
            when "10" & x"7d6" => DATA <= x"fa8f";
            when "10" & x"7d7" => DATA <= x"a8ff";
            when "10" & x"7d8" => DATA <= x"805f";
            when "10" & x"7d9" => DATA <= x"e032";
            when "10" & x"7da" => DATA <= x"0984";
            when "10" & x"7db" => DATA <= x"0744";
            when "10" & x"7dc" => DATA <= x"0000";
            when "10" & x"7dd" => DATA <= x"1c80";
            when "10" & x"7de" => DATA <= x"2058";
            when "10" & x"7df" => DATA <= x"0807";
            when "10" & x"7e0" => DATA <= x"4181";
            when "10" & x"7e1" => DATA <= x"d55c";
            when "10" & x"7e2" => DATA <= x"15fe";
            when "10" & x"7e3" => DATA <= x"dd7f";
            when "10" & x"7e4" => DATA <= x"c8fb";
            when "10" & x"7e5" => DATA <= x"f0c6";
            when "10" & x"7e6" => DATA <= x"7c7e";
            when "10" & x"7e7" => DATA <= x"1888";
            when "10" & x"7e8" => DATA <= x"0f87";
            when "10" & x"7e9" => DATA <= x"e3f5";
            when "10" & x"7ea" => DATA <= x"3efd";
            when "10" & x"7eb" => DATA <= x"7a9f";
            when "10" & x"7ec" => DATA <= x"4f67";
            when "10" & x"7ed" => DATA <= x"93d1";
            when "10" & x"7ee" => DATA <= x"fc92";
            when "10" & x"7ef" => DATA <= x"0200";
            when "10" & x"7f0" => DATA <= x"b800";
            when "10" & x"7f1" => DATA <= x"00a3";
            when "10" & x"7f2" => DATA <= x"2480";
            when "10" & x"7f3" => DATA <= x"3fc0";
            when "10" & x"7f4" => DATA <= x"0424";
            when "10" & x"7f5" => DATA <= x"6180";
            when "10" & x"7f6" => DATA <= x"f048";
            when "10" & x"7f7" => DATA <= x"383f";
            when "10" & x"7f8" => DATA <= x"e800";
            when "10" & x"7f9" => DATA <= x"6067";
            when "10" & x"7fa" => DATA <= x"141e";
            when "10" & x"7fb" => DATA <= x"0dcf";
            when "10" & x"7fc" => DATA <= x"b023";
            when "10" & x"7fd" => DATA <= x"8c00";
            when "10" & x"7fe" => DATA <= x"02ac";
            when "10" & x"7ff" => DATA <= x"0700";
            when "10" & x"800" => DATA <= x"fc21";
            when "10" & x"801" => DATA <= x"4000";
            when "10" & x"802" => DATA <= x"e7f8";
            when "10" & x"803" => DATA <= x"0680";
            when "10" & x"804" => DATA <= x"0094";
            when "10" & x"805" => DATA <= x"0050";
            when "10" & x"806" => DATA <= x"7fa1";
            when "10" & x"807" => DATA <= x"9001";
            when "10" & x"808" => DATA <= x"0507";
            when "10" & x"809" => DATA <= x"003f";
            when "10" & x"80a" => DATA <= x"c007";
            when "10" & x"80b" => DATA <= x"f280";
            when "10" & x"80c" => DATA <= x"8000";
            when "10" & x"80d" => DATA <= x"8000";
            when "10" & x"80e" => DATA <= x"35c6";
            when "10" & x"80f" => DATA <= x"00f0";
            when "10" & x"810" => DATA <= x"39c0";
            when "10" & x"811" => DATA <= x"0007";
            when "10" & x"812" => DATA <= x"003f";
            when "10" & x"813" => DATA <= x"c80c";
            when "10" & x"814" => DATA <= x"6703";
            when "10" & x"815" => DATA <= x"89c8";
            when "10" & x"816" => DATA <= x"cc00";
            when "10" & x"817" => DATA <= x"1fda";
            when "10" & x"818" => DATA <= x"93fe";
            when "10" & x"819" => DATA <= x"2400";
            when "10" & x"81a" => DATA <= x"3fcf";
            when "10" & x"81b" => DATA <= x"f3fe";
            when "10" & x"81c" => DATA <= x"fc00";
            when "10" & x"81d" => DATA <= x"3fe8";
            when "10" & x"81e" => DATA <= x"0106";
            when "10" & x"81f" => DATA <= x"8700";
            when "10" & x"820" => DATA <= x"2000";
            when "10" & x"821" => DATA <= x"00ba";
            when "10" & x"822" => DATA <= x"0040";
            when "10" & x"823" => DATA <= x"2601";
            when "10" & x"824" => DATA <= x"0297";
            when "10" & x"825" => DATA <= x"f006";
            when "10" & x"826" => DATA <= x"8000";
            when "10" & x"827" => DATA <= x"6fda";
            when "10" & x"828" => DATA <= x"027f";
            when "10" & x"829" => DATA <= x"c803";
            when "10" & x"82a" => DATA <= x"fe80";
            when "10" & x"82b" => DATA <= x"1ff2";
            when "10" & x"82c" => DATA <= x"00ff";
            when "10" & x"82d" => DATA <= x"a017";
            when "10" & x"82e" => DATA <= x"fd78";
            when "10" & x"82f" => DATA <= x"1e11";
            when "10" & x"830" => DATA <= x"0ffa";
            when "10" & x"831" => DATA <= x"00af";
            when "10" & x"832" => DATA <= x"f3f9";
            when "10" & x"833" => DATA <= x"584a";
            when "10" & x"834" => DATA <= x"ff00";
            when "10" & x"835" => DATA <= x"081f";
            when "10" & x"836" => DATA <= x"f5fc";
            when "10" & x"837" => DATA <= x"004f";
            when "10" & x"838" => DATA <= x"bfc0";
            when "10" & x"839" => DATA <= x"0f37";
            when "10" & x"83a" => DATA <= x"f804";
            when "10" & x"83b" => DATA <= x"febe";
            when "10" & x"83c" => DATA <= x"aff1";
            when "10" & x"83d" => DATA <= x"c009";
            when "10" & x"83e" => DATA <= x"fe00";
            when "10" & x"83f" => DATA <= x"013f";
            when "10" & x"840" => DATA <= x"12a5";
            when "10" & x"841" => DATA <= x"f020";
            when "10" & x"842" => DATA <= x"01ff";
            when "10" & x"843" => DATA <= x"400f";
            when "10" & x"844" => DATA <= x"f571";
            when "10" & x"845" => DATA <= x"f000";
            when "10" & x"846" => DATA <= x"20a0";
            when "10" & x"847" => DATA <= x"05c3";
            when "10" & x"848" => DATA <= x"e402";
            when "10" & x"849" => DATA <= x"c700";
            when "10" & x"84a" => DATA <= x"011e";
            when "10" & x"84b" => DATA <= x"000a";
            when "10" & x"84c" => DATA <= x"ff70";
            when "10" & x"84d" => DATA <= x"2140";
            when "10" & x"84e" => DATA <= x"4007";
            when "10" & x"84f" => DATA <= x"f801";
            when "10" & x"850" => DATA <= x"f6bf";
            when "10" & x"851" => DATA <= x"7780";
            when "10" & x"852" => DATA <= x"1f40";
            when "10" & x"853" => DATA <= x"07f8";
            when "10" & x"854" => DATA <= x"01fa";
            when "10" & x"855" => DATA <= x"257f";
            when "10" & x"856" => DATA <= x"be9f";
            when "10" & x"857" => DATA <= x"ee03";
            when "10" & x"858" => DATA <= x"f800";
            when "10" & x"859" => DATA <= x"7ef1";
            when "10" & x"85a" => DATA <= x"7f87";
            when "10" & x"85b" => DATA <= x"cfe8";
            when "10" & x"85c" => DATA <= x"7e00";
            when "10" & x"85d" => DATA <= x"0e93";
            when "10" & x"85e" => DATA <= x"df8e";
            when "10" & x"85f" => DATA <= x"6707";
            when "10" & x"860" => DATA <= x"0007";
            when "10" & x"861" => DATA <= x"2c02";
            when "10" & x"862" => DATA <= x"8200";
            when "10" & x"863" => DATA <= x"0f87";
            when "10" & x"864" => DATA <= x"8006";
            when "10" & x"865" => DATA <= x"802b";
            when "10" & x"866" => DATA <= x"f800";
            when "10" & x"867" => DATA <= x"dc20";
            when "10" & x"868" => DATA <= x"2728";
            when "10" & x"869" => DATA <= x"01fe";
            when "10" & x"86a" => DATA <= x"fe00";
            when "10" & x"86b" => DATA <= x"3cde";
            when "10" & x"86c" => DATA <= x"2020";
            when "10" & x"86d" => DATA <= x"0311";
            when "10" & x"86e" => DATA <= x"8e07";
            when "10" & x"86f" => DATA <= x"000f";
            when "10" & x"870" => DATA <= x"c394";
            when "10" & x"871" => DATA <= x"0001";
            when "10" & x"872" => DATA <= x"3fd2";
            when "10" & x"873" => DATA <= x"0107";
            when "10" & x"874" => DATA <= x"8005";
            when "10" & x"875" => DATA <= x"1400";
            when "10" & x"876" => DATA <= x"40a0";
            when "10" & x"877" => DATA <= x"0010";
            when "10" & x"878" => DATA <= x"0007";
            when "10" & x"879" => DATA <= x"6002";
            when "10" & x"87a" => DATA <= x"0030";
            when "10" & x"87b" => DATA <= x"0020";
            when "10" & x"87c" => DATA <= x"0078";
            when "10" & x"87d" => DATA <= x"5002";
            when "10" & x"87e" => DATA <= x"4e40";
            when "10" & x"87f" => DATA <= x"1ce8";
            when "10" & x"880" => DATA <= x"2400";
            when "10" & x"881" => DATA <= x"0801";
            when "10" & x"882" => DATA <= x"4020";
            when "10" & x"883" => DATA <= x"2758";
            when "10" & x"884" => DATA <= x"0004";
            when "10" & x"885" => DATA <= x"4000";
            when "10" & x"886" => DATA <= x"1028";
            when "10" & x"887" => DATA <= x"008d";
            when "10" & x"888" => DATA <= x"4000";
            when "10" & x"889" => DATA <= x"1900";
            when "10" & x"88a" => DATA <= x"7ad0";
            when "10" & x"88b" => DATA <= x"02c2";
            when "10" & x"88c" => DATA <= x"b010";
            when "10" & x"88d" => DATA <= x"0887";
            when "10" & x"88e" => DATA <= x"7001";
            when "10" & x"88f" => DATA <= x"e002";
            when "10" & x"890" => DATA <= x"9000";
            when "10" & x"891" => DATA <= x"0998";
            when "10" & x"892" => DATA <= x"00fe";
            when "10" & x"893" => DATA <= x"7ccf";
            when "10" & x"894" => DATA <= x"f9fc";
            when "10" & x"895" => DATA <= x"f150";
            when "10" & x"896" => DATA <= x"7c06";
            when "10" & x"897" => DATA <= x"4341";
            when "10" & x"898" => DATA <= x"80c7";
            when "10" & x"899" => DATA <= x"e079";
            when "10" & x"89a" => DATA <= x"000c";
            when "10" & x"89b" => DATA <= x"1f9e";
            when "10" & x"89c" => DATA <= x"0720";
            when "10" & x"89d" => DATA <= x"5020";
            when "10" & x"89e" => DATA <= x"0006";
            when "10" & x"89f" => DATA <= x"7082";
            when "10" & x"8a0" => DATA <= x"0072";
            when "10" & x"8a1" => DATA <= x"0080";
            when "10" & x"8a2" => DATA <= x"0688";
            when "10" & x"8a3" => DATA <= x"2c1d";
            when "10" & x"8a4" => DATA <= x"7ef7";
            when "10" & x"8a5" => DATA <= x"7803";
            when "10" & x"8a6" => DATA <= x"2b12";
            when "10" & x"8a7" => DATA <= x"8017";
            when "10" & x"8a8" => DATA <= x"d5fe";
            when "10" & x"8a9" => DATA <= x"2423";
            when "10" & x"8aa" => DATA <= x"31a8";
            when "10" & x"8ab" => DATA <= x"016d";
            when "10" & x"8ac" => DATA <= x"5fe0";
            when "10" & x"8ad" => DATA <= x"2001";
            when "10" & x"8ae" => DATA <= x"9a80";
            when "10" & x"8af" => DATA <= x"1ed5";
            when "10" & x"8b0" => DATA <= x"fe00";
            when "10" & x"8b1" => DATA <= x"5f70";
            when "10" & x"8b2" => DATA <= x"03d9";
            when "10" & x"8b3" => DATA <= x"febf";
            when "10" & x"8b4" => DATA <= x"0020";
            when "10" & x"8b5" => DATA <= x"d08a";
            when "10" & x"8b6" => DATA <= x"0003";
            when "10" & x"8b7" => DATA <= x"b9de";
            when "10" & x"8b8" => DATA <= x"3308";
            when "10" & x"8b9" => DATA <= x"0480";
            when "10" & x"8ba" => DATA <= x"9c00";
            when "10" & x"8bb" => DATA <= x"0770";
            when "10" & x"8bc" => DATA <= x"5003";
            when "10" & x"8bd" => DATA <= x"9a80";
            when "10" & x"8be" => DATA <= x"0404";
            when "10" & x"8bf" => DATA <= x"0140";
            when "10" & x"8c0" => DATA <= x"2012";
            when "10" & x"8c1" => DATA <= x"6801";
            when "10" & x"8c2" => DATA <= x"1298";
            when "10" & x"8c3" => DATA <= x"0004";
            when "10" & x"8c4" => DATA <= x"7a05";
            when "10" & x"8c5" => DATA <= x"fe77";
            when "10" & x"8c6" => DATA <= x"42bd";
            when "10" & x"8c7" => DATA <= x"c060";
            when "10" & x"8c8" => DATA <= x"0240";
            when "10" & x"8c9" => DATA <= x"201e";
            when "10" & x"8ca" => DATA <= x"4231";
            when "10" & x"8cb" => DATA <= x"bfce";
            when "10" & x"8cc" => DATA <= x"0000";
            when "10" & x"8cd" => DATA <= x"c380";
            when "10" & x"8ce" => DATA <= x"0046";
            when "10" & x"8cf" => DATA <= x"603f";
            when "10" & x"8d0" => DATA <= x"db80";
            when "10" & x"8d1" => DATA <= x"0402";
            when "10" & x"8d2" => DATA <= x"4dbe";
            when "10" & x"8d3" => DATA <= x"8c44";
            when "10" & x"8d4" => DATA <= x"2244";
            when "10" & x"8d5" => DATA <= x"2807";
            when "10" & x"8d6" => DATA <= x"9b0e";
            when "10" & x"8d7" => DATA <= x"bc07";
            when "10" & x"8d8" => DATA <= x"03f4";
            when "10" & x"8d9" => DATA <= x"181d";
            when "10" & x"8da" => DATA <= x"40b0";
            when "10" & x"8db" => DATA <= x"0198";
            when "10" & x"8dc" => DATA <= x"1402";
            when "10" & x"8dd" => DATA <= x"407b";
            when "10" & x"8de" => DATA <= x"91f0";
            when "10" & x"8df" => DATA <= x"f0ef";
            when "10" & x"8e0" => DATA <= x"87eb";
            when "10" & x"8e1" => DATA <= x"f1fe";
            when "10" & x"8e2" => DATA <= x"c723";
            when "10" & x"8e3" => DATA <= x"81c0";
            when "10" & x"8e4" => DATA <= x"607e";
            when "10" & x"8e5" => DATA <= x"0300";
            when "10" & x"8e6" => DATA <= x"a02b";
            when "10" & x"8e7" => DATA <= x"fa40";
            when "10" & x"8e8" => DATA <= x"11d5";
            when "10" & x"8e9" => DATA <= x"1e81";
            when "10" & x"8ea" => DATA <= x"a80a";
            when "10" & x"8eb" => DATA <= x"00fd";
            when "10" & x"8ec" => DATA <= x"f7fd";
            when "10" & x"8ed" => DATA <= x"fb85";
            when "10" & x"8ee" => DATA <= x"c032";
            when "10" & x"8ef" => DATA <= x"e340";
            when "10" & x"8f0" => DATA <= x"2000";
            when "10" & x"8f1" => DATA <= x"0d0e";
            when "10" & x"8f2" => DATA <= x"0783";
            when "10" & x"8f3" => DATA <= x"9c00";
            when "10" & x"8f4" => DATA <= x"1cde";
            when "10" & x"8f5" => DATA <= x"f000";
            when "10" & x"8f6" => DATA <= x"0ddf";
            when "10" & x"8f7" => DATA <= x"47d4";
            when "10" & x"8f8" => DATA <= x"3c3e";
            when "10" & x"8f9" => DATA <= x"a001";
            when "10" & x"8fa" => DATA <= x"f006";
            when "10" & x"8fb" => DATA <= x"4007";
            when "10" & x"8fc" => DATA <= x"880a";
            when "10" & x"8fd" => DATA <= x"0040";
            when "10" & x"8fe" => DATA <= x"4803";
            when "10" & x"8ff" => DATA <= x"fde0";
            when "10" & x"900" => DATA <= x"c0ae";
            when "10" & x"901" => DATA <= x"0525";
            when "10" & x"902" => DATA <= x"7257";
            when "10" & x"903" => DATA <= x"3a74";
            when "10" & x"904" => DATA <= x"3e5f";
            when "10" & x"905" => DATA <= x"2f17";
            when "10" & x"906" => DATA <= x"c3e9";
            when "10" & x"907" => DATA <= x"f0eb";
            when "10" & x"908" => DATA <= x"b240";
            when "10" & x"909" => DATA <= x"2a00";
            when "10" & x"90a" => DATA <= x"00fa";
            when "10" & x"90b" => DATA <= x"72b8";
            when "10" & x"90c" => DATA <= x"1f8f";
            when "10" & x"90d" => DATA <= x"77a3";
            when "10" & x"90e" => DATA <= x"d5e8";
            when "10" & x"90f" => DATA <= x"b640";
            when "10" & x"910" => DATA <= x"8041";
            when "10" & x"911" => DATA <= x"a150";
            when "10" & x"912" => DATA <= x"2820";
            when "10" & x"913" => DATA <= x"0081";
            when "10" & x"914" => DATA <= x"420a";
            when "10" & x"915" => DATA <= x"0005";
            when "10" & x"916" => DATA <= x"4e00";
            when "10" & x"917" => DATA <= x"0108";
            when "10" & x"918" => DATA <= x"8920";
            when "10" & x"919" => DATA <= x"0380";
            when "10" & x"91a" => DATA <= x"0426";
            when "10" & x"91b" => DATA <= x"8804";
            when "10" & x"91c" => DATA <= x"0415";
            when "10" & x"91d" => DATA <= x"6002";
            when "10" & x"91e" => DATA <= x"bd00";
            when "10" & x"91f" => DATA <= x"1802";
            when "10" & x"920" => DATA <= x"0002";
            when "10" & x"921" => DATA <= x"e240";
            when "10" & x"922" => DATA <= x"d140";
            when "10" & x"923" => DATA <= x"00ca";
            when "10" & x"924" => DATA <= x"004a";
            when "10" & x"925" => DATA <= x"0107";
            when "10" & x"926" => DATA <= x"cc0a";
            when "10" & x"927" => DATA <= x"0060";
            when "10" & x"928" => DATA <= x"2016";
            when "10" & x"929" => DATA <= x"a006";
            when "10" & x"92a" => DATA <= x"6001";
            when "10" & x"92b" => DATA <= x"2010";
            when "10" & x"92c" => DATA <= x"a000";
            when "10" & x"92d" => DATA <= x"9001";
            when "10" & x"92e" => DATA <= x"bfc0";
            when "10" & x"92f" => DATA <= x"0c03";
            when "10" & x"930" => DATA <= x"0300";
            when "10" & x"931" => DATA <= x"0038";
            when "10" & x"932" => DATA <= x"0051";
            when "10" & x"933" => DATA <= x"0190";
            when "10" & x"934" => DATA <= x"88ff";
            when "10" & x"935" => DATA <= x"0004";
            when "10" & x"936" => DATA <= x"7800";
            when "10" & x"937" => DATA <= x"02f0";
            when "10" & x"938" => DATA <= x"6d00";
            when "10" & x"939" => DATA <= x"0ae0";
            when "10" & x"93a" => DATA <= x"0a80";
            when "10" & x"93b" => DATA <= x"0018";
            when "10" & x"93c" => DATA <= x"4e02";
            when "10" & x"93d" => DATA <= x"05e8";
            when "10" & x"93e" => DATA <= x"0008";
            when "10" & x"93f" => DATA <= x"0040";
            when "10" & x"940" => DATA <= x"29c7";
            when "10" & x"941" => DATA <= x"2134";
            when "10" & x"942" => DATA <= x"7700";
            when "10" & x"943" => DATA <= x"220b";
            when "10" & x"944" => DATA <= x"a3f0";
            when "10" & x"945" => DATA <= x"0958";
            when "10" & x"946" => DATA <= x"0011";
            when "10" & x"947" => DATA <= x"a030";
            when "10" & x"948" => DATA <= x"1101";
            when "10" & x"949" => DATA <= x"8200";
            when "10" & x"94a" => DATA <= x"0870";
            when "10" & x"94b" => DATA <= x"075e";
            when "10" & x"94c" => DATA <= x"bf45";
            when "10" & x"94d" => DATA <= x"0240";
            when "10" & x"94e" => DATA <= x"20a1";
            when "10" & x"94f" => DATA <= x"ccc0";
            when "10" & x"950" => DATA <= x"64bb";
            when "10" & x"951" => DATA <= x"cc34";
            when "10" & x"952" => DATA <= x"0010";
            when "10" & x"953" => DATA <= x"2000";
            when "10" & x"954" => DATA <= x"02e0";
            when "10" & x"955" => DATA <= x"1033";
            when "10" & x"956" => DATA <= x"e190";
            when "10" & x"957" => DATA <= x"a80f";
            when "10" & x"958" => DATA <= x"4800";
            when "10" & x"959" => DATA <= x"5002";
            when "10" & x"95a" => DATA <= x"c003";
            when "10" & x"95b" => DATA <= x"b808";
            when "10" & x"95c" => DATA <= x"0100";
            when "10" & x"95d" => DATA <= x"037c";
            when "10" & x"95e" => DATA <= x"0080";
            when "10" & x"95f" => DATA <= x"00a0";
            when "10" & x"960" => DATA <= x"530f";
            when "10" & x"961" => DATA <= x"c002";
            when "10" & x"962" => DATA <= x"fb80";
            when "10" & x"963" => DATA <= x"17c9";
            when "10" & x"964" => DATA <= x"a578";
            when "10" & x"965" => DATA <= x"017e";
            when "10" & x"966" => DATA <= x"3038";
            when "10" & x"967" => DATA <= x"021b";
            when "10" & x"968" => DATA <= x"0fd7";
            when "10" & x"969" => DATA <= x"f00c";
            when "10" & x"96a" => DATA <= x"3c80";
            when "10" & x"96b" => DATA <= x"a000";
            when "10" & x"96c" => DATA <= x"081d";
            when "10" & x"96d" => DATA <= x"6090";
            when "10" & x"96e" => DATA <= x"0800";
            when "10" & x"96f" => DATA <= x"6400";
            when "10" & x"970" => DATA <= x"220f";
            when "10" & x"971" => DATA <= x"d000";
            when "10" & x"972" => DATA <= x"1018";
            when "10" & x"973" => DATA <= x"0404";
            when "10" & x"974" => DATA <= x"063e";
            when "10" & x"975" => DATA <= x"2800";
            when "10" & x"976" => DATA <= x"c000";
            when "10" & x"977" => DATA <= x"7850";
            when "10" & x"978" => DATA <= x"03fc";
            when "10" & x"979" => DATA <= x"1c10";
            when "10" & x"97a" => DATA <= x"0250";
            when "10" & x"97b" => DATA <= x"0260";
            when "10" & x"97c" => DATA <= x"61dc";
            when "10" & x"97d" => DATA <= x"6fc7";
            when "10" & x"97e" => DATA <= x"8b82";
            when "10" & x"97f" => DATA <= x"8018";
            when "10" & x"980" => DATA <= x"1440";
            when "10" & x"981" => DATA <= x"0804";
            when "10" & x"982" => DATA <= x"bbc0";
            when "10" & x"983" => DATA <= x"0200";
            when "10" & x"984" => DATA <= x"0801";
            when "10" & x"985" => DATA <= x"0000";
            when "10" & x"986" => DATA <= x"4005";
            when "10" & x"987" => DATA <= x"c03c";
            when "10" & x"988" => DATA <= x"0088";
            when "10" & x"989" => DATA <= x"403e";
            when "10" & x"98a" => DATA <= x"000c";
            when "10" & x"98b" => DATA <= x"0407";
            when "10" & x"98c" => DATA <= x"241b";
            when "10" & x"98d" => DATA <= x"9fe3";
            when "10" & x"98e" => DATA <= x"2020";
            when "10" & x"98f" => DATA <= x"0002";
            when "10" & x"990" => DATA <= x"2108";
            when "10" & x"991" => DATA <= x"001f";
            when "10" & x"992" => DATA <= x"e0ee";
            when "10" & x"993" => DATA <= x"0023";
            when "10" & x"994" => DATA <= x"9201";
            when "10" & x"995" => DATA <= x"0ff0";
            when "10" & x"996" => DATA <= x"0024";
            when "10" & x"997" => DATA <= x"07c1";
            when "10" & x"998" => DATA <= x"00a0";
            when "10" & x"999" => DATA <= x"0a82";
            when "10" & x"99a" => DATA <= x"8014";
            when "10" & x"99b" => DATA <= x"1400";
            when "10" & x"99c" => DATA <= x"c000";
            when "10" & x"99d" => DATA <= x"0044";
            when "10" & x"99e" => DATA <= x"c042";
            when "10" & x"99f" => DATA <= x"1d00";
            when "10" & x"9a0" => DATA <= x"3fe4";
            when "10" & x"9a1" => DATA <= x"0025";
            when "10" & x"9a2" => DATA <= x"200c";
            when "10" & x"9a3" => DATA <= x"0240";
            when "10" & x"9a4" => DATA <= x"2000";
            when "10" & x"9a5" => DATA <= x"0ee0";
            when "10" & x"9a6" => DATA <= x"01a5";
            when "10" & x"9a7" => DATA <= x"0010";
            when "10" & x"9a8" => DATA <= x"827c";
            when "10" & x"9a9" => DATA <= x"007d";
            when "10" & x"9aa" => DATA <= x"580c";
            when "10" & x"9ab" => DATA <= x"000d";
            when "10" & x"9ac" => DATA <= x"5125";
            when "10" & x"9ad" => DATA <= x"0032";
            when "10" & x"9ae" => DATA <= x"4008";
            when "10" & x"9af" => DATA <= x"0623";
            when "10" & x"9b0" => DATA <= x"7f80";
            when "10" & x"9b1" => DATA <= x"1c4e";
            when "10" & x"9b2" => DATA <= x"061b";
            when "10" & x"9b3" => DATA <= x"f501";
            when "10" & x"9b4" => DATA <= x"c01c";
            when "10" & x"9b5" => DATA <= x"3eff";
            when "10" & x"9b6" => DATA <= x"7cd7";
            when "10" & x"9b7" => DATA <= x"c578";
            when "10" & x"9b8" => DATA <= x"3e1e";
            when "10" & x"9b9" => DATA <= x"0231";
            when "10" & x"9ba" => DATA <= x"ef0e";
            when "10" & x"9bb" => DATA <= x"80c5";
            when "10" & x"9bc" => DATA <= x"609f";
            when "10" & x"9bd" => DATA <= x"00a0";
            when "10" & x"9be" => DATA <= x"0024";
            when "10" & x"9bf" => DATA <= x"8001";
            when "10" & x"9c0" => DATA <= x"3c02";
            when "10" & x"9c1" => DATA <= x"803c";
            when "10" & x"9c2" => DATA <= x"1c0e";
            when "10" & x"9c3" => DATA <= x"0e27";
            when "10" & x"9c4" => DATA <= x"0780";
            when "10" & x"9c5" => DATA <= x"406a";
            when "10" & x"9c6" => DATA <= x"0e05";
            when "10" & x"9c7" => DATA <= x"7805";
            when "10" & x"9c8" => DATA <= x"0051";
            when "10" & x"9c9" => DATA <= x"4500";
            when "10" & x"9ca" => DATA <= x"0a94";
            when "10" & x"9cb" => DATA <= x"1c00";
            when "10" & x"9cc" => DATA <= x"42a0";
            when "10" & x"9cd" => DATA <= x"0204";
            when "10" & x"9ce" => DATA <= x"8004";
            when "10" & x"9cf" => DATA <= x"2800";
            when "10" & x"9d0" => DATA <= x"2140";
            when "10" & x"9d1" => DATA <= x"0040";
            when "10" & x"9d2" => DATA <= x"6012";
            when "10" & x"9d3" => DATA <= x"8300";
            when "10" & x"9d4" => DATA <= x"9419";
            when "10" & x"9d5" => DATA <= x"e000";
            when "10" & x"9d6" => DATA <= x"0b01";
            when "10" & x"9d7" => DATA <= x"0180";
            when "10" & x"9d8" => DATA <= x"6800";
            when "10" & x"9d9" => DATA <= x"83c0";
            when "10" & x"9da" => DATA <= x"010e";
            when "10" & x"9db" => DATA <= x"0000";
            when "10" & x"9dc" => DATA <= x"e801";
            when "10" & x"9dd" => DATA <= x"8000";
            when "10" & x"9de" => DATA <= x"02e0";
            when "10" & x"9df" => DATA <= x"0040";
            when "10" & x"9e0" => DATA <= x"0103";
            when "10" & x"9e1" => DATA <= x"a00c";
            when "10" & x"9e2" => DATA <= x"0005";
            when "10" & x"9e3" => DATA <= x"71bf";
            when "10" & x"9e4" => DATA <= x"dde8";
            when "10" & x"9e5" => DATA <= x"f7fa";
            when "10" & x"9e6" => DATA <= x"7dfe";
            when "10" & x"9e7" => DATA <= x"ef37";
            when "10" & x"9e8" => DATA <= x"bbdf";
            when "10" & x"9e9" => DATA <= x"e0f3";
            when "10" & x"9ea" => DATA <= x"7950";
            when "10" & x"9eb" => DATA <= x"6ef8";
            when "10" & x"9ec" => DATA <= x"7c8c";
            when "10" & x"9ed" => DATA <= x"9f13";
            when "10" & x"9ee" => DATA <= x"f340";
            when "10" & x"9ef" => DATA <= x"7586";
            when "10" & x"9f0" => DATA <= x"c7a0";
            when "10" & x"9f1" => DATA <= x"303b";
            when "10" & x"9f2" => DATA <= x"edfc";
            when "10" & x"9f3" => DATA <= x"ff07";
            when "10" & x"9f4" => DATA <= x"8058";
            when "10" & x"9f5" => DATA <= x"15fc";
            when "10" & x"9f6" => DATA <= x"9200";
            when "10" & x"9f7" => DATA <= x"80d0";
            when "10" & x"9f8" => DATA <= x"08e4";
            when "10" & x"9f9" => DATA <= x"7a1d";
            when "10" & x"9fa" => DATA <= x"0007";
            when "10" & x"9fb" => DATA <= x"0030";
            when "10" & x"9fc" => DATA <= x"377c";
            when "10" & x"9fd" => DATA <= x"00f0";
            when "10" & x"9fe" => DATA <= x"bf70";
            when "10" & x"9ff" => DATA <= x"0146";
            when "10" & x"a00" => DATA <= x"dc43";
            when "10" & x"a01" => DATA <= x"943c";
            when "10" & x"a02" => DATA <= x"1c0f";
            when "10" & x"a03" => DATA <= x"70e3";
            when "10" & x"a04" => DATA <= x"bebf";
            when "10" & x"a05" => DATA <= x"f7bc";
            when "10" & x"a06" => DATA <= x"7d47";
            when "10" & x"a07" => DATA <= x"fa7c";
            when "10" & x"a08" => DATA <= x"1f7f";
            when "10" & x"a09" => DATA <= x"f00a";
            when "10" & x"a0a" => DATA <= x"e280";
            when "10" & x"a0b" => DATA <= x"4c00";
            when "10" & x"a0c" => DATA <= x"3e00";
            when "10" & x"a0d" => DATA <= x"66d0";
            when "10" & x"a0e" => DATA <= x"0570";
            when "10" & x"a0f" => DATA <= x"301c";
            when "10" & x"a10" => DATA <= x"0804";
            when "10" & x"a11" => DATA <= x"ea01";
            when "10" & x"a12" => DATA <= x"c123";
            when "10" & x"a13" => DATA <= x"e1b0";
            when "10" & x"a14" => DATA <= x"fb6d";
            when "10" & x"a15" => DATA <= x"be00";
            when "10" & x"a16" => DATA <= x"4000";
            when "10" & x"a17" => DATA <= x"008d";
            when "10" & x"a18" => DATA <= x"4edc";
            when "10" & x"a19" => DATA <= x"7fbd";
            when "10" & x"a1a" => DATA <= x"3bf1";
            when "10" & x"a1b" => DATA <= x"faf4";
            when "10" & x"a1c" => DATA <= x"7a81";
            when "10" & x"a1d" => DATA <= x"000f";
            when "10" & x"a1e" => DATA <= x"f017";
            when "10" & x"a1f" => DATA <= x"0180";
            when "10" & x"a20" => DATA <= x"0040";
            when "10" & x"a21" => DATA <= x"073b";
            when "10" & x"a22" => DATA <= x"c2c0";
            when "10" & x"a23" => DATA <= x"1fa0";
            when "10" & x"a24" => DATA <= x"5a04";
            when "10" & x"a25" => DATA <= x"0101";
            when "10" & x"a26" => DATA <= x"00c0";
            when "10" & x"a27" => DATA <= x"01b9";
            when "10" & x"a28" => DATA <= x"02c0";
            when "10" & x"a29" => DATA <= x"17e1";
            when "10" & x"a2a" => DATA <= x"ba08";
            when "10" & x"a2b" => DATA <= x"0270";
            when "10" & x"a2c" => DATA <= x"013d";
            when "10" & x"a2d" => DATA <= x"0160";
            when "10" & x"a2e" => DATA <= x"0ee1";
            when "10" & x"a2f" => DATA <= x"7d10";
            when "10" & x"a30" => DATA <= x"0404";
            when "10" & x"a31" => DATA <= x"0300";
            when "10" & x"a32" => DATA <= x"02fc";
            when "10" & x"a33" => DATA <= x"0022";
            when "10" & x"a34" => DATA <= x"0008";
            when "10" & x"a35" => DATA <= x"3801";
            when "10" & x"a36" => DATA <= x"b8da";
            when "10" & x"a37" => DATA <= x"2110";
            when "10" & x"a38" => DATA <= x"045c";
            when "10" & x"a39" => DATA <= x"007d";
            when "10" & x"a3a" => DATA <= x"f003";
            when "10" & x"a3b" => DATA <= x"d892";
            when "10" & x"a3c" => DATA <= x"8010";
            when "10" & x"a3d" => DATA <= x"0004";
            when "10" & x"a3e" => DATA <= x"0001";
            when "10" & x"a3f" => DATA <= x"efc0";
            when "10" & x"a40" => DATA <= x"2000";
            when "10" & x"a41" => DATA <= x"0d00";
            when "10" & x"a42" => DATA <= x"3d5a";
            when "10" & x"a43" => DATA <= x"1400";
            when "10" & x"a44" => DATA <= x"11e0";
            when "10" & x"a45" => DATA <= x"07f8";
            when "10" & x"a46" => DATA <= x"1a80";
            when "10" & x"a47" => DATA <= x"8020";
            when "10" & x"a48" => DATA <= x"0010";
            when "10" & x"a49" => DATA <= x"0136";
            when "10" & x"a4a" => DATA <= x"e0b0";
            when "10" & x"a4b" => DATA <= x"07d8";
            when "10" & x"a4c" => DATA <= x"2682";
            when "10" & x"a4d" => DATA <= x"0080";
            when "10" & x"a4e" => DATA <= x"8020";
            when "10" & x"a4f" => DATA <= x"005e";
            when "10" & x"a50" => DATA <= x"c0b0";
            when "10" & x"a51" => DATA <= x"07b8";
            when "10" & x"a52" => DATA <= x"5a84";
            when "10" & x"a53" => DATA <= x"1d01";
            when "10" & x"a54" => DATA <= x"000a";
            when "10" & x"a55" => DATA <= x"a002";
            when "10" & x"a56" => DATA <= x"0701";
            when "10" & x"a57" => DATA <= x"0000";
            when "10" & x"a58" => DATA <= x"2000";
            when "10" & x"a59" => DATA <= x"8060";
            when "10" & x"a5a" => DATA <= x"07c0";
            when "10" & x"a5b" => DATA <= x"0ff1";
            when "10" & x"a5c" => DATA <= x"cd80";
            when "10" & x"a5d" => DATA <= x"3fc0";
            when "10" & x"a5e" => DATA <= x"4007";
            when "10" & x"a5f" => DATA <= x"09e4";
            when "10" & x"a60" => DATA <= x"5143";
            when "10" & x"a61" => DATA <= x"0732";
            when "10" & x"a62" => DATA <= x"61c0";
            when "10" & x"a63" => DATA <= x"e280";
            when "10" & x"a64" => DATA <= x"380c";
            when "10" & x"a65" => DATA <= x"0e0f";
            when "10" & x"a66" => DATA <= x"0e00";
            when "10" & x"a67" => DATA <= x"7ff0";
            when "10" & x"a68" => DATA <= x"200c";
            when "10" & x"a69" => DATA <= x"0802";
            when "10" & x"a6a" => DATA <= x"0025";
            when "10" & x"a6b" => DATA <= x"c814";
            when "10" & x"a6c" => DATA <= x"0040";
            when "10" & x"a6d" => DATA <= x"e005";
            when "10" & x"a6e" => DATA <= x"d86e";
            when "10" & x"a6f" => DATA <= x"8200";
            when "10" & x"a70" => DATA <= x"808a";
            when "10" & x"a71" => DATA <= x"0027";
            when "10" & x"a72" => DATA <= x"a02c";
            when "10" & x"a73" => DATA <= x"01dc";
            when "10" & x"a74" => DATA <= x"2fa2";
            when "10" & x"a75" => DATA <= x"0080";
            when "10" & x"a76" => DATA <= x"0060";
            when "10" & x"a77" => DATA <= x"007f";
            when "10" & x"a78" => DATA <= x"d801";
            when "10" & x"a79" => DATA <= x"01f8";
            when "10" & x"a7a" => DATA <= x"dba4";
            when "10" & x"a7b" => DATA <= x"0101";
            when "10" & x"a7c" => DATA <= x"0280";
            when "10" & x"a7d" => DATA <= x"0fbe";
            when "10" & x"a7e" => DATA <= x"00f3";
            when "10" & x"a7f" => DATA <= x"5a50";
            when "10" & x"a80" => DATA <= x"0200";
            when "10" & x"a81" => DATA <= x"0080";
            when "10" & x"a82" => DATA <= x"003f";
            when "10" & x"a83" => DATA <= x"f806";
            when "10" & x"a84" => DATA <= x"8000";
            when "10" & x"a85" => DATA <= x"2007";
            when "10" & x"a86" => DATA <= x"2b62";
            when "10" & x"a87" => DATA <= x"c01f";
            when "10" & x"a88" => DATA <= x"fc04";
            when "10" & x"a89" => DATA <= x"0501";
            when "10" & x"a8a" => DATA <= x"0040";
            when "10" & x"a8b" => DATA <= x"0fb5";
            when "10" & x"a8c" => DATA <= x"0580";
            when "10" & x"a8d" => DATA <= x"36c1";
            when "10" & x"a8e" => DATA <= x"b410";
            when "10" & x"a8f" => DATA <= x"04e0";
            when "10" & x"a90" => DATA <= x"01f9";
            when "10" & x"a91" => DATA <= x"02c0";
            when "10" & x"a92" => DATA <= x"1ee1";
            when "10" & x"a93" => DATA <= x"6a10";
            when "10" & x"a94" => DATA <= x"0404";
            when "10" & x"a95" => DATA <= x"0300";
            when "10" & x"a96" => DATA <= x"06ff";
            when "10" & x"a97" => DATA <= x"803f";
            when "10" & x"a98" => DATA <= x"cdb4";
            when "10" & x"a99" => DATA <= x"4120";
            when "10" & x"a9a" => DATA <= x"0ffd";
            when "10" & x"a9b" => DATA <= x"0006";
            when "10" & x"a9c" => DATA <= x"0017";
            when "10" & x"a9d" => DATA <= x"3501";
            when "10" & x"a9e" => DATA <= x"4008";
            when "10" & x"a9f" => DATA <= x"04f0";
            when "10" & x"aa0" => DATA <= x"7bbf";
            when "10" & x"aa1" => DATA <= x"a9f8";
            when "10" & x"aa2" => DATA <= x"eaf0";
            when "10" & x"aa3" => DATA <= x"7f1f";
            when "10" & x"aa4" => DATA <= x"c1e0";
            when "10" & x"aa5" => DATA <= x"1e00";
            when "10" & x"aa6" => DATA <= x"a69a";
            when "10" & x"aa7" => DATA <= x"0834";
            when "10" & x"aa8" => DATA <= x"0200";
            when "10" & x"aa9" => DATA <= x"030f";
            when "10" & x"aaa" => DATA <= x"0000";
            when "10" & x"aab" => DATA <= x"5025";
            when "10" & x"aac" => DATA <= x"0001";
            when "10" & x"aad" => DATA <= x"3801";
            when "10" & x"aae" => DATA <= x"81c0";
            when "10" & x"aaf" => DATA <= x"040e";
            when "10" & x"ab0" => DATA <= x"0007";
            when "10" & x"ab1" => DATA <= x"f839";
            when "10" & x"ab2" => DATA <= x"203d";
            when "10" & x"ab3" => DATA <= x"41c0";
            when "10" & x"ab4" => DATA <= x"a0f5";
            when "10" & x"ab5" => DATA <= x"0778";
            when "10" & x"ab6" => DATA <= x"0000";
            when "10" & x"ab7" => DATA <= x"54aa";
            when "10" & x"ab8" => DATA <= x"0008";
            when "10" & x"ab9" => DATA <= x"000a";
            when "10" & x"aba" => DATA <= x"8a00";
            when "10" & x"abb" => DATA <= x"2006";
            when "10" & x"abc" => DATA <= x"3800";
            when "10" & x"abd" => DATA <= x"8140";
            when "10" & x"abe" => DATA <= x"0140";
            when "10" & x"abf" => DATA <= x"8700";
            when "10" & x"ac0" => DATA <= x"0428";
            when "10" & x"ac1" => DATA <= x"000d";
            when "10" & x"ac2" => DATA <= x"4180";
            when "10" & x"ac3" => DATA <= x"4a0c";
            when "10" & x"ac4" => DATA <= x"0203";
            when "10" & x"ac5" => DATA <= x"3c00";
            when "10" & x"ac6" => DATA <= x"0140";
            when "10" & x"ac7" => DATA <= x"203d";
            when "10" & x"ac8" => DATA <= x"0128";
            when "10" & x"ac9" => DATA <= x"7000";
            when "10" & x"aca" => DATA <= x"07c0";
            when "10" & x"acb" => DATA <= x"2400";
            when "10" & x"acc" => DATA <= x"0540";
            when "10" & x"acd" => DATA <= x"0081";
            when "10" & x"ace" => DATA <= x"1680";
            when "10" & x"acf" => DATA <= x"2024";
            when "10" & x"ad0" => DATA <= x"0101";
            when "10" & x"ad1" => DATA <= x"5fe9";
            when "10" & x"ad2" => DATA <= x"f7ff";
            when "10" & x"ad3" => DATA <= x"6fa7";
            when "10" & x"ad4" => DATA <= x"def4";
            when "10" & x"ad5" => DATA <= x"2fbe";
            when "10" & x"ad6" => DATA <= x"ef6a";
            when "10" & x"ad7" => DATA <= x"ff7f";
            when "10" & x"ad8" => DATA <= x"3e1b";
            when "10" & x"ad9" => DATA <= x"0187";
            when "10" & x"ada" => DATA <= x"c681";
            when "10" & x"adb" => DATA <= x"d61b";
            when "10" & x"adc" => DATA <= x"1e40";
            when "10" & x"add" => DATA <= x"1fcf";
            when "10" & x"ade" => DATA <= x"f078";
            when "10" & x"adf" => DATA <= x"0100";
            when "10" & x"ae0" => DATA <= x"00a8";
            when "10" & x"ae1" => DATA <= x"0408";
            when "10" & x"ae2" => DATA <= x"0c00";
            when "10" & x"ae3" => DATA <= x"8cad";
            when "10" & x"ae4" => DATA <= x"faff";
            when "10" & x"ae5" => DATA <= x"0180";
            when "10" & x"ae6" => DATA <= x"1a0d";
            when "10" & x"ae7" => DATA <= x"faf7";
            when "10" & x"ae8" => DATA <= x"7f80";
            when "10" & x"ae9" => DATA <= x"d800";
            when "10" & x"aea" => DATA <= x"0af7";
            when "10" & x"aeb" => DATA <= x"38d0";
            when "10" & x"aec" => DATA <= x"0800";
            when "10" & x"aed" => DATA <= x"0200";
            when "10" & x"aee" => DATA <= x"009c";
            when "10" & x"aef" => DATA <= x"7800";
            when "10" & x"af0" => DATA <= x"3c1c";
            when "10" & x"af1" => DATA <= x"e1e7";
            when "10" & x"af2" => DATA <= x"7d00";
            when "10" & x"af3" => DATA <= x"3beb";
            when "10" & x"af4" => DATA <= x"febb";
            when "10" & x"af5" => DATA <= x"c7d4";
            when "10" & x"af6" => DATA <= x"01c7";
            when "10" & x"af7" => DATA <= x"e3e0";
            when "10" & x"af8" => DATA <= x"f005";
            when "10" & x"af9" => DATA <= x"8000";
            when "10" & x"afa" => DATA <= x"1e3f";
            when "10" & x"afb" => DATA <= x"2401";
            when "10" & x"afc" => DATA <= x"fe70";
            when "10" & x"afd" => DATA <= x"4003";
            when "10" & x"afe" => DATA <= x"f801";
            when "10" & x"aff" => DATA <= x"815c";
            when "10" & x"b00" => DATA <= x"0e77";
            when "10" & x"b01" => DATA <= x"3572";
            when "10" & x"b02" => DATA <= x"292b";
            when "10" & x"b03" => DATA <= x"7c3e";
            when "10" & x"b04" => DATA <= x"dde1";
            when "10" & x"b05" => DATA <= x"f4f5";
            when "10" & x"b06" => DATA <= x"7a3f";
            when "10" & x"b07" => DATA <= x"2a70";
            when "10" & x"b08" => DATA <= x"2815";
            when "10" & x"b09" => DATA <= x"4a3f";
            when "10" & x"b0a" => DATA <= x"5ecf";
            when "10" & x"b0b" => DATA <= x"faf7";
            when "10" & x"b0c" => DATA <= x"7ed7";
            when "10" & x"b0d" => DATA <= x"ff80";
            when "10" & x"b0e" => DATA <= x"7804";
            when "10" & x"b0f" => DATA <= x"8050";
            when "10" & x"b10" => DATA <= x"2002";
            when "10" & x"b11" => DATA <= x"813c";
            when "10" & x"b12" => DATA <= x"03c0";
            when "10" & x"b13" => DATA <= x"3c02";
            when "10" & x"b14" => DATA <= x"c004";
            when "10" & x"b15" => DATA <= x"1401";
            when "10" & x"b16" => DATA <= x"441e";
            when "10" & x"b17" => DATA <= x"01e0";
            when "10" & x"b18" => DATA <= x"1e01";
            when "10" & x"b19" => DATA <= x"e01e";
            when "10" & x"b1a" => DATA <= x"01c0";
            when "10" & x"b1b" => DATA <= x"001f";
            when "10" & x"b1c" => DATA <= x"00f0";
            when "10" & x"b1d" => DATA <= x"0f00";
            when "10" & x"b1e" => DATA <= x"f000";
            when "10" & x"b1f" => DATA <= x"4780";
            when "10" & x"b20" => DATA <= x"7800";
            when "10" & x"b21" => DATA <= x"0021";
            when "10" & x"b22" => DATA <= x"4001";
            when "10" & x"b23" => DATA <= x"0b00";
            when "10" & x"b24" => DATA <= x"0470";
            when "10" & x"b25" => DATA <= x"0064";
            when "10" & x"b26" => DATA <= x"6239";
            when "10" & x"b27" => DATA <= x"04d1";
            when "10" & x"b28" => DATA <= x"c864";
            when "10" & x"b29" => DATA <= x"3b20";
            when "10" & x"b2a" => DATA <= x"040e";
            when "10" & x"b2b" => DATA <= x"0022";
            when "10" & x"b2c" => DATA <= x"5269";
            when "10" & x"b2d" => DATA <= x"1293";
            when "10" & x"b2e" => DATA <= x"4884";
            when "10" & x"b2f" => DATA <= x"df00";
            when "10" & x"b30" => DATA <= x"f00f";
            when "10" & x"b31" => DATA <= x"00f0";
            when "10" & x"b32" => DATA <= x"0000";
            when "10" & x"b33" => DATA <= x"23c0";
            when "10" & x"b34" => DATA <= x"3400";
            when "10" & x"b35" => DATA <= x"4140";
            when "10" & x"b36" => DATA <= x"020f";
            when "10" & x"b37" => DATA <= x"00f0";
            when "10" & x"b38" => DATA <= x"0001";
            when "10" & x"b39" => DATA <= x"03c0";
            when "10" & x"b3a" => DATA <= x"3c03";
            when "10" & x"b3b" => DATA <= x"c03c";
            when "10" & x"b3c" => DATA <= x"03c0";
            when "10" & x"b3d" => DATA <= x"0000";
            when "10" & x"b3e" => DATA <= x"2a00";
            when "10" & x"b3f" => DATA <= x"0178";
            when "10" & x"b40" => DATA <= x"0780";
            when "10" & x"b41" => DATA <= x"7807";
            when "10" & x"b42" => DATA <= x"8004";
            when "10" & x"b43" => DATA <= x"2802";
            when "10" & x"b44" => DATA <= x"843c";
            when "10" & x"b45" => DATA <= x"03c0";
            when "10" & x"b46" => DATA <= x"3c02";
            when "10" & x"b47" => DATA <= x"403e";
            when "10" & x"b48" => DATA <= x"0101";
            when "10" & x"b49" => DATA <= x"2f94";
            when "10" & x"b4a" => DATA <= x"fa7c";
            when "10" & x"b4b" => DATA <= x"3ed6";
            when "10" & x"b4c" => DATA <= x"03e1";
            when "10" & x"b4d" => DATA <= x"b0f8";
            when "10" & x"b4e" => DATA <= x"7857";
            when "10" & x"b4f" => DATA <= x"c06c";
            when "10" & x"b50" => DATA <= x"f743";
            when "10" & x"b51" => DATA <= x"74f6";
            when "10" & x"b52" => DATA <= x"1b1d";
            when "10" & x"b53" => DATA <= x"f805";
            when "10" & x"b54" => DATA <= x"0001";
            when "10" & x"b55" => DATA <= x"2802";
            when "10" & x"b56" => DATA <= x"8100";
            when "10" & x"b57" => DATA <= x"0040";
            when "10" & x"b58" => DATA <= x"0103";
            when "10" & x"b59" => DATA <= x"8008";
            when "10" & x"b5a" => DATA <= x"1400";
            when "10" & x"b5b" => DATA <= x"0707";
            when "10" & x"b5c" => DATA <= x"f038";
            when "10" & x"b5d" => DATA <= x"3e81";
            when "10" & x"b5e" => DATA <= x"c1d4";
            when "10" & x"b5f" => DATA <= x"0002";
            when "10" & x"b60" => DATA <= x"2f10";
            when "10" & x"b61" => DATA <= x"0040";
            when "10" & x"b62" => DATA <= x"ef00";
            when "10" & x"b63" => DATA <= x"008a";
            when "10" & x"b64" => DATA <= x"a801";
            when "10" & x"b65" => DATA <= x"4028";
            when "10" & x"b66" => DATA <= x"5500";
            when "10" & x"b67" => DATA <= x"1504";
            when "10" & x"b68" => DATA <= x"0e00";
            when "10" & x"b69" => DATA <= x"a400";
            when "10" & x"b6a" => DATA <= x"0100";
            when "10" & x"b6b" => DATA <= x"ab40";
            when "10" & x"b6c" => DATA <= x"0140";
            when "10" & x"b6d" => DATA <= x"8054";
            when "10" & x"b6e" => DATA <= x"0054";
            when "10" & x"b6f" => DATA <= x"0203";
            when "10" & x"b70" => DATA <= x"b830";
            when "10" & x"b71" => DATA <= x"1c04";
            when "10" & x"b72" => DATA <= x"0670";
            when "10" & x"b73" => DATA <= x"0202";
            when "10" & x"b74" => DATA <= x"4028";
            when "10" & x"b75" => DATA <= x"0400";
            when "10" & x"b76" => DATA <= x"03a0";
            when "10" & x"b77" => DATA <= x"1005";
            when "10" & x"b78" => DATA <= x"0080";
            when "10" & x"b79" => DATA <= x"0025";
            when "10" & x"b7a" => DATA <= x"4a00";
            when "10" & x"b7b" => DATA <= x"0080";
            when "10" & x"b7c" => DATA <= x"0020";
            when "10" & x"b7d" => DATA <= x"000a";
            when "10" & x"b7e" => DATA <= x"8280";
            when "10" & x"b7f" => DATA <= x"0020";
            when "10" & x"b80" => DATA <= x"0510";
            when "10" & x"b81" => DATA <= x"0104";
            when "10" & x"b82" => DATA <= x"2a10";
            when "10" & x"b83" => DATA <= x"0000";
            when "10" & x"b84" => DATA <= x"4000";
            when "10" & x"b85" => DATA <= x"8000";
            when "10" & x"b86" => DATA <= x"20c0";
            when "10" & x"b87" => DATA <= x"a000";
            when "10" & x"b88" => DATA <= x"8203";
            when "10" & x"b89" => DATA <= x"8fc3";
            when "10" & x"b8a" => DATA <= x"f47e";
            when "10" & x"b8b" => DATA <= x"bf4f";
            when "10" & x"b8c" => DATA <= x"810e";
            when "10" & x"b8d" => DATA <= x"e040";
            when "10" & x"b8e" => DATA <= x"ba5c";
            when "10" & x"b8f" => DATA <= x"2cc5";
            when "10" & x"b90" => DATA <= x"47be";
            when "10" & x"b91" => DATA <= x"5f0f";
            when "10" & x"b92" => DATA <= x"9048";
            when "10" & x"b93" => DATA <= x"1dfc";
            when "10" & x"b94" => DATA <= x"ff3f";
            when "10" & x"b95" => DATA <= x"80d8";
            when "10" & x"b96" => DATA <= x"740e";
            when "10" & x"b97" => DATA <= x"4001";
            when "10" & x"b98" => DATA <= x"81c4";
            when "10" & x"b99" => DATA <= x"0c07";
            when "10" & x"b9a" => DATA <= x"fbf9";
            when "10" & x"b9b" => DATA <= x"bc00";
            when "10" & x"b9c" => DATA <= x"0230";
            when "10" & x"b9d" => DATA <= x"1c15";
            when "10" & x"b9e" => DATA <= x"1e81";
            when "10" & x"b9f" => DATA <= x"4900";
            when "10" & x"ba0" => DATA <= x"100f";
            when "10" & x"ba1" => DATA <= x"77fe";
            when "10" & x"ba2" => DATA <= x"efbf";
            when "10" & x"ba3" => DATA <= x"d40f";
            when "10" & x"ba4" => DATA <= x"fdf7";
            when "10" & x"ba5" => DATA <= x"7f80";
            when "10" & x"ba6" => DATA <= x"1fe7";
            when "10" & x"ba7" => DATA <= x"118c";
            when "10" & x"ba8" => DATA <= x"b89c";
            when "10" & x"ba9" => DATA <= x"0e34";
            when "10" & x"baa" => DATA <= x"3d43";
            when "10" & x"bab" => DATA <= x"9c00";
            when "10" & x"bac" => DATA <= x"1e9e";
            when "10" & x"bad" => DATA <= x"fa00";
            when "10" & x"bae" => DATA <= x"77bf";
            when "10" & x"baf" => DATA <= x"d3c1";
            when "10" & x"bb0" => DATA <= x"ea3e";
            when "10" & x"bb1" => DATA <= x"a001";
            when "10" & x"bb2" => DATA <= x"f0fc";
            when "10" & x"bb3" => DATA <= x"77c0";
            when "10" & x"bb4" => DATA <= x"0f80";
            when "10" & x"bb5" => DATA <= x"003d";
            when "10" & x"bb6" => DATA <= x"feef";
            when "10" & x"bb7" => DATA <= x"e007";
            when "10" & x"bb8" => DATA <= x"fbc0";
            when "10" & x"bb9" => DATA <= x"8007";
            when "10" & x"bba" => DATA <= x"7629";
            when "10" & x"bbb" => DATA <= x"2b92";
            when "10" & x"bbc" => DATA <= x"b9dc";
            when "10" & x"bbd" => DATA <= x"0f00";
            when "10" & x"bbe" => DATA <= x"fa78";
            when "10" & x"bbf" => DATA <= x"3e9f";
            when "10" & x"bc0" => DATA <= x"0f87";
            when "10" & x"bc1" => DATA <= x"13e1";
            when "10" & x"bc2" => DATA <= x"f4a2";
            when "10" & x"bc3" => DATA <= x"543a";
            when "10" & x"bc4" => DATA <= x"15a9";
            when "10" & x"bc5" => DATA <= x"448a";
            when "10" & x"bc6" => DATA <= x"51fe";
            when "10" & x"bc7" => DATA <= x"fdaf";
            when "10" & x"bc8" => DATA <= x"f7a3";
            when "10" & x"bc9" => DATA <= x"c1ea";
            when "10" & x"bca" => DATA <= x"f490";
            when "10" & x"bcb" => DATA <= x"0187";
            when "10" & x"bcc" => DATA <= x"8020";
            when "10" & x"bcd" => DATA <= x"3800";
            when "10" & x"bce" => DATA <= x"09a0";
            when "10" & x"bcf" => DATA <= x"004f";
            when "10" & x"bd0" => DATA <= x"00f0";
            when "10" & x"bd1" => DATA <= x"0f00";
            when "10" & x"bd2" => DATA <= x"9001";
            when "10" & x"bd3" => DATA <= x"0680";
            when "10" & x"bd4" => DATA <= x"0834";
            when "10" & x"bd5" => DATA <= x"0005";
            when "10" & x"bd6" => DATA <= x"e000";
            when "10" & x"bd7" => DATA <= x"8f00";
            when "10" & x"bd8" => DATA <= x"f00f";
            when "10" & x"bd9" => DATA <= x"00f0";
            when "10" & x"bda" => DATA <= x"0e00";
            when "10" & x"bdb" => DATA <= x"2078";
            when "10" & x"bdc" => DATA <= x"0043";
            when "10" & x"bdd" => DATA <= x"c03c";
            when "10" & x"bde" => DATA <= x"0380";
            when "10" & x"bdf" => DATA <= x"011e";
            when "10" & x"be0" => DATA <= x"01e0";
            when "10" & x"be1" => DATA <= x"0000";
            when "10" & x"be2" => DATA <= x"8780";
            when "10" & x"be3" => DATA <= x"5000";
            when "10" & x"be4" => DATA <= x"26a6";
            when "10" & x"be5" => DATA <= x"4320";
            when "10" & x"be6" => DATA <= x"1a39";
            when "10" & x"be7" => DATA <= x"04d8";
            when "10" & x"be8" => DATA <= x"0008";
            when "10" & x"be9" => DATA <= x"0045";
            when "10" & x"bea" => DATA <= x"a4c2";
            when "10" & x"beb" => DATA <= x"6902";
            when "10" & x"bec" => DATA <= x"9348";
            when "10" & x"bed" => DATA <= x"9200";
            when "10" & x"bee" => DATA <= x"0ff0";
            when "10" & x"bef" => DATA <= x"0a00";
            when "10" & x"bf0" => DATA <= x"0278";
            when "10" & x"bf1" => DATA <= x"0500";
            when "10" & x"bf2" => DATA <= x"5045";
            when "10" & x"bf3" => DATA <= x"0006";
            when "10" & x"bf4" => DATA <= x"3c03";
            when "10" & x"bf5" => DATA <= x"c000";
            when "10" & x"bf6" => DATA <= x"030f";
            when "10" & x"bf7" => DATA <= x"00f0";
            when "10" & x"bf8" => DATA <= x"0003";
            when "10" & x"bf9" => DATA <= x"0000";
            when "10" & x"bfa" => DATA <= x"40f0";
            when "10" & x"bfb" => DATA <= x"0b00";
            when "10" & x"bfc" => DATA <= x"4078";
            when "10" & x"bfd" => DATA <= x"0007";
            when "10" & x"bfe" => DATA <= x"c024";
            when "10" & x"bff" => DATA <= x"0280";
            when "10" & x"c00" => DATA <= x"a800";
            when "10" & x"c01" => DATA <= x"0c00";
            when "10" & x"c02" => DATA <= x"0178";
            when "10" & x"c03" => DATA <= x"0580";
            when "10" & x"c04" => DATA <= x"033c";
            when "10" & x"c05" => DATA <= x"0240";
            when "10" & x"c06" => DATA <= x"021c";
            when "10" & x"c07" => DATA <= x"0038";
            when "10" & x"c08" => DATA <= x"0004";
            when "10" & x"c09" => DATA <= x"3c02";
            when "10" & x"c0a" => DATA <= x"c00c";
            when "10" & x"c0b" => DATA <= x"1e01";
            when "10" & x"c0c" => DATA <= x"201f";
            when "10" & x"c0d" => DATA <= x"0080";
            when "10" & x"c0e" => DATA <= x"3e9f";
            when "10" & x"c0f" => DATA <= x"0e9c";
            when "10" & x"c10" => DATA <= x"f94f";
            when "10" & x"c11" => DATA <= x"b5f1";
            when "10" & x"c12" => DATA <= x"5b15";
            when "10" & x"c13" => DATA <= x"f0f0";
            when "10" & x"c14" => DATA <= x"6c50";
            when "10" & x"c15" => DATA <= x"d82c";
            when "10" & x"c16" => DATA <= x"363b";
            when "10" & x"c17" => DATA <= x"159a";
            when "10" & x"c18" => DATA <= x"c77e";
            when "10" & x"c19" => DATA <= x"01a0";
            when "10" & x"c1a" => DATA <= x"0040";
            when "10" & x"c1b" => DATA <= x"0502";
            when "10" & x"c1c" => DATA <= x"5801";
            when "10" & x"c1d" => DATA <= x"0001";
            when "10" & x"c1e" => DATA <= x"60e0";
            when "10" & x"c1f" => DATA <= x"f33e";
            when "10" & x"c20" => DATA <= x"8000";
            when "10" & x"c21" => DATA <= x"881e";
            when "10" & x"c22" => DATA <= x"0140";
            when "10" & x"c23" => DATA <= x"0a0a";
            when "10" & x"c24" => DATA <= x"0040";
            when "10" & x"c25" => DATA <= x"5000";
            when "10" & x"c26" => DATA <= x"a800";
            when "10" & x"c27" => DATA <= x"40b0";
            when "10" & x"c28" => DATA <= x"0200";
            when "10" & x"c29" => DATA <= x"1280";
            when "10" & x"c2a" => DATA <= x"0034";
            when "10" & x"c2b" => DATA <= x"0015";
            when "10" & x"c2c" => DATA <= x"0081";
            when "10" & x"c2d" => DATA <= x"3430";
            when "10" & x"c2e" => DATA <= x"0c0c";
            when "10" & x"c2f" => DATA <= x"f00a";
            when "10" & x"c30" => DATA <= x"00a0";
            when "10" & x"c31" => DATA <= x"1000";
            when "10" & x"c32" => DATA <= x"0f80";
            when "10" & x"c33" => DATA <= x"6800";
            when "10" & x"c34" => DATA <= x"2140";
            when "10" & x"c35" => DATA <= x"010f";
            when "10" & x"c36" => DATA <= x"0000";
            when "10" & x"c37" => DATA <= x"0068";
            when "10" & x"c38" => DATA <= x"0050";
            when "10" & x"c39" => DATA <= x"0ae0";
            when "10" & x"c3a" => DATA <= x"0547";
            when "10" & x"c3b" => DATA <= x"0004";
            when "10" & x"c3c" => DATA <= x"000c";
            when "10" & x"c3d" => DATA <= x"0000";
            when "10" & x"c3e" => DATA <= x"4100";
            when "10" & x"c3f" => DATA <= x"9f5f";
            when "10" & x"c40" => DATA <= x"a7d7";
            when "10" & x"c41" => DATA <= x"e9fa";
            when "10" & x"c42" => DATA <= x"bf4f";
            when "10" & x"c43" => DATA <= x"ab74";
            when "10" & x"c44" => DATA <= x"b43a";
            when "10" & x"c45" => DATA <= x"9d7f";
            when "10" & x"c46" => DATA <= x"9f0f";
            when "10" & x"c47" => DATA <= x"d2f8";
            when "10" & x"c48" => DATA <= x"fca0";
            when "10" & x"c49" => DATA <= x"07c2";
            when "10" & x"c4a" => DATA <= x"2801";
            when "10" & x"c4b" => DATA <= x"4201";
            when "10" & x"c4c" => DATA <= x"37ab";
            when "10" & x"c4d" => DATA <= x"3008";
            when "10" & x"c4e" => DATA <= x"3400";
            when "10" & x"c4f" => DATA <= x"1fce";
            when "10" & x"c50" => DATA <= x"47fa";
            when "10" & x"c51" => DATA <= x"ff7e";
            when "10" & x"c52" => DATA <= x"6ff7";
            when "10" & x"c53" => DATA <= x"ffff";
            when "10" & x"c54" => DATA <= x"fd7f";
            when "10" & x"c55" => DATA <= x"d388";
            when "10" & x"c56" => DATA <= x"c75c";
            when "10" & x"c57" => DATA <= x"43d4";
            when "10" & x"c58" => DATA <= x"381e";
            when "10" & x"c59" => DATA <= x"a1ca";
            when "10" & x"c5a" => DATA <= x"1eff";
            when "10" & x"c5b" => DATA <= x"f7fc";
            when "10" & x"c5c" => DATA <= x"9fcf";
            when "10" & x"c5d" => DATA <= x"ff00";
            when "10" & x"c5e" => DATA <= x"bf00";
            when "10" & x"c5f" => DATA <= x"6010";
            when "10" & x"c60" => DATA <= x"0083";
            when "10" & x"c61" => DATA <= x"801f";
            when "10" & x"c62" => DATA <= x"e800";
            when "10" & x"c63" => DATA <= x"2098";
            when "10" & x"c64" => DATA <= x"18c0";
            when "10" & x"c65" => DATA <= x"7020";
            when "10" & x"c66" => DATA <= x"13b3";
            when "10" & x"c67" => DATA <= x"815b";
            when "10" & x"c68" => DATA <= x"edb0";
            when "10" & x"c69" => DATA <= x"fa7f";
            when "10" & x"c6a" => DATA <= x"87da";
            when "10" & x"c6b" => DATA <= x"89c6";
            when "10" & x"c6c" => DATA <= x"a362";
            when "10" & x"c6d" => DATA <= x"b41e";
            when "10" & x"c6e" => DATA <= x"8d4f";
            when "10" & x"c6f" => DATA <= x"f77a";
            when "10" & x"c70" => DATA <= x"f807";
            when "10" & x"c71" => DATA <= x"8070";
            when "10" & x"c72" => DATA <= x"0502";
            when "10" & x"c73" => DATA <= x"0000";
            when "10" & x"c74" => DATA <= x"9400";
            when "10" & x"c75" => DATA <= x"04f0";
            when "10" & x"c76" => DATA <= x"0f00";
            when "10" & x"c77" => DATA <= x"f009";
            when "10" & x"c78" => DATA <= x"0010";
            when "10" & x"c79" => DATA <= x"5005";
            when "10" & x"c7a" => DATA <= x"1000";
            when "10" & x"c7b" => DATA <= x"041e";
            when "10" & x"c7c" => DATA <= x"01e0";
            when "10" & x"c7d" => DATA <= x"1e01";
            when "10" & x"c7e" => DATA <= x"e01e";
            when "10" & x"c7f" => DATA <= x"01e0";
            when "10" & x"c80" => DATA <= x"1e01";
            when "10" & x"c81" => DATA <= x"e01e";
            when "10" & x"c82" => DATA <= x"01e0";
            when "10" & x"c83" => DATA <= x"1e01";
            when "10" & x"c84" => DATA <= x"2001";
            when "10" & x"c85" => DATA <= x"0f00";
            when "10" & x"c86" => DATA <= x"f00a";
            when "10" & x"c87" => DATA <= x"3900";
            when "10" & x"c88" => DATA <= x"8e68";
            when "10" & x"c89" => DATA <= x"6472";
            when "10" & x"c8a" => DATA <= x"0900";
            when "10" & x"c8b" => DATA <= x"1000";
            when "10" & x"c8c" => DATA <= x"0029";
            when "10" & x"c8d" => DATA <= x"0026";
            when "10" & x"c8e" => DATA <= x"9308";
            when "10" & x"c8f" => DATA <= x"84c2";
            when "10" & x"c90" => DATA <= x"6f26";
            when "10" & x"c91" => DATA <= x"7805";
            when "10" & x"c92" => DATA <= x"0001";
            when "10" & x"c93" => DATA <= x"3c03";
            when "10" & x"c94" => DATA <= x"c03c";
            when "10" & x"c95" => DATA <= x"03c0";
            when "10" & x"c96" => DATA <= x"3c03";
            when "10" & x"c97" => DATA <= x"c03c";
            when "10" & x"c98" => DATA <= x"0000";
            when "10" & x"c99" => DATA <= x"40f0";
            when "10" & x"c9a" => DATA <= x"0f00";
            when "10" & x"c9b" => DATA <= x"f00f";
            when "10" & x"c9c" => DATA <= x"00f0";
            when "10" & x"c9d" => DATA <= x"0000";
            when "10" & x"c9e" => DATA <= x"0b40";
            when "10" & x"c9f" => DATA <= x"005e";
            when "10" & x"ca0" => DATA <= x"01e0";
            when "10" & x"ca1" => DATA <= x"1e01";
            when "10" & x"ca2" => DATA <= x"2001";
            when "10" & x"ca3" => DATA <= x"0e00";
            when "10" & x"ca4" => DATA <= x"0878";
            when "10" & x"ca5" => DATA <= x"0780";
            when "10" & x"ca6" => DATA <= x"7806";
            when "10" & x"ca7" => DATA <= x"807c";
            when "10" & x"ca8" => DATA <= x"0200";
            when "10" & x"ca9" => DATA <= x"fa1c";
            when "10" & x"caa" => DATA <= x"2e0f";
            when "10" & x"cab" => DATA <= x"5faf";
            when "10" & x"cac" => DATA <= x"c7eb";
            when "10" & x"cad" => DATA <= x"7420";
            when "10" & x"cae" => DATA <= x"60a0";
            when "10" & x"caf" => DATA <= x"0a01";
            when "10" & x"cb0" => DATA <= x"0401";
            when "10" & x"cb1" => DATA <= x"0343";
            when "10" & x"cb2" => DATA <= x"a181";
            when "10" & x"cb3" => DATA <= x"61f0";
            when "10" & x"cb4" => DATA <= x"002a";
            when "10" & x"cb5" => DATA <= x"4803";
            when "10" & x"cb6" => DATA <= x"3d7e";
            when "10" & x"cb7" => DATA <= x"005e";
            when "10" & x"cb8" => DATA <= x"c803";
            when "10" & x"cb9" => DATA <= x"fc62";
            when "10" & x"cba" => DATA <= x"307d";
            when "10" & x"cbb" => DATA <= x"c801";
            when "10" & x"cbc" => DATA <= x"e400";
            when "10" & x"cbd" => DATA <= x"701e";
            when "10" & x"cbe" => DATA <= x"8100";
            when "10" & x"cbf" => DATA <= x"e470";
            when "10" & x"cc0" => DATA <= x"387c";
            when "10" & x"cc1" => DATA <= x"1f43";
            when "10" & x"cc2" => DATA <= x"e3ff";
            when "10" & x"cc3" => DATA <= x"0028";
            when "10" & x"cc4" => DATA <= x"7804";
            when "10" & x"cc5" => DATA <= x"802a";
            when "10" & x"cc6" => DATA <= x"3800";
            when "10" & x"cc7" => DATA <= x"41c0";
            when "10" & x"cc8" => DATA <= x"042e";
            when "10" & x"cc9" => DATA <= x"0020";
            when "10" & x"cca" => DATA <= x"7001";
            when "10" & x"ccb" => DATA <= x"5000";
            when "10" & x"ccc" => DATA <= x"01a0";
            when "10" & x"ccd" => DATA <= x"0060";
            when "10" & x"cce" => DATA <= x"1283";
            when "10" & x"ccf" => DATA <= x"0080";
            when "10" & x"cd0" => DATA <= x"c020";
            when "10" & x"cd1" => DATA <= x"33c0";
            when "10" & x"cd2" => DATA <= x"0012";
            when "10" & x"cd3" => DATA <= x"0200";
            when "10" & x"cd4" => DATA <= x"e01a";
            when "10" & x"cd5" => DATA <= x"0000";
            when "10" & x"cd6" => DATA <= x"8000";
            when "10" & x"cd7" => DATA <= x"3a00";
            when "10" & x"cd8" => DATA <= x"a1d0";
            when "10" & x"cd9" => DATA <= x"0045";
            when "10" & x"cda" => DATA <= x"0170";
            when "10" & x"cdb" => DATA <= x"0008";
            when "10" & x"cdc" => DATA <= x"0080";
            when "10" & x"cdd" => DATA <= x"0004";
            when "10" & x"cde" => DATA <= x"2801";
            when "10" & x"cdf" => DATA <= x"0140";
            when "10" & x"ce0" => DATA <= x"01fe";
            when "10" & x"ce1" => DATA <= x"3f07";
            when "10" & x"ce2" => DATA <= x"b9eb";
            when "10" & x"ce3" => DATA <= x"3d3a";
            when "10" & x"ce4" => DATA <= x"9b4f";
            when "10" & x"ce5" => DATA <= x"83d1";
            when "10" & x"ce6" => DATA <= x"ead7";
            when "10" & x"ce7" => DATA <= x"0a04";
            when "10" & x"ce8" => DATA <= x"01df";
            when "10" & x"ce9" => DATA <= x"94fe";
            when "10" & x"cea" => DATA <= x"5f3f";
            when "10" & x"ceb" => DATA <= x"a028";
            when "10" & x"cec" => DATA <= x"0ce7";
            when "10" & x"ced" => DATA <= x"2009";
            when "10" & x"cee" => DATA <= x"6693";
            when "10" & x"cef" => DATA <= x"696c";
            when "10" & x"cf0" => DATA <= x"0400";
            when "10" & x"cf1" => DATA <= x"57e3";
            when "10" & x"cf2" => DATA <= x"fdf0";
            when "10" & x"cf3" => DATA <= x"fa7d";
            when "10" & x"cf4" => DATA <= x"a000";
            when "10" & x"cf5" => DATA <= x"0850";
            when "10" & x"cf6" => DATA <= x"1dff";
            when "10" & x"cf7" => DATA <= x"83c0";
            when "10" & x"cf8" => DATA <= x"1bfe";
            when "10" & x"cf9" => DATA <= x"0768";
            when "10" & x"cfa" => DATA <= x"0029";
            when "10" & x"cfb" => DATA <= x"c4a3";
            when "10" & x"cfc" => DATA <= x"4020";
            when "10" & x"cfd" => DATA <= x"0008";
            when "10" & x"cfe" => DATA <= x"0287";
            when "10" & x"cff" => DATA <= x"b872";
            when "10" & x"d00" => DATA <= x"8783";
            when "10" & x"d01" => DATA <= x"9fff";
            when "10" & x"d02" => DATA <= x"bff4";
            when "10" & x"d03" => DATA <= x"7f57";
            when "10" & x"d04" => DATA <= x"e210";
            when "10" & x"d05" => DATA <= x"3d00";
            when "10" & x"d06" => DATA <= x"f003";
            when "10" & x"d07" => DATA <= x"fe82";
            when "10" & x"d08" => DATA <= x"150e";
            when "10" & x"d09" => DATA <= x"8e00";
            when "10" & x"d0a" => DATA <= x"7fd6";
            when "10" & x"d0b" => DATA <= x"033d";
            when "10" & x"d0c" => DATA <= x"8ce4";
            when "10" & x"d0d" => DATA <= x"6138";
            when "10" & x"d0e" => DATA <= x"1812";
            when "10" & x"d0f" => DATA <= x"3e9f";
            when "10" & x"d10" => DATA <= x"a1f0";
            when "10" & x"d11" => DATA <= x"f341";
            when "10" & x"d12" => DATA <= x"295a";
            when "10" & x"d13" => DATA <= x"0d56";
            when "10" & x"d14" => DATA <= x"2d6a";
            when "10" & x"d15" => DATA <= x"3dfb";
            when "10" & x"d16" => DATA <= x"d5ee";
            when "10" & x"d17" => DATA <= x"f5af";
            when "10" & x"d18" => DATA <= x"7f00";
            when "10" & x"d19" => DATA <= x"f00a";
            when "10" & x"d1a" => DATA <= x"0002";
            when "10" & x"d1b" => DATA <= x"5000";
            when "10" & x"d1c" => DATA <= x"1380";
            when "10" & x"d1d" => DATA <= x"009e";
            when "10" & x"d1e" => DATA <= x"01e0";
            when "10" & x"d1f" => DATA <= x"1e01";
            when "10" & x"d20" => DATA <= x"c002";
            when "10" & x"d21" => DATA <= x"0a00";
            when "10" & x"d22" => DATA <= x"1000";
            when "10" & x"d23" => DATA <= x"0400";
            when "10" & x"d24" => DATA <= x"0107";
            when "10" & x"d25" => DATA <= x"8078";
            when "10" & x"d26" => DATA <= x"0780";
            when "10" & x"d27" => DATA <= x"7807";
            when "10" & x"d28" => DATA <= x"8078";
            when "10" & x"d29" => DATA <= x"0580";
            when "10" & x"d2a" => DATA <= x"00bc";
            when "10" & x"d2b" => DATA <= x"03c0";
            when "10" & x"d2c" => DATA <= x"2400";
            when "10" & x"d2d" => DATA <= x"11e0";
            when "10" & x"d2e" => DATA <= x"1e00";
            when "10" & x"d2f" => DATA <= x"0008";
            when "10" & x"d30" => DATA <= x"7800";
            when "10" & x"d31" => DATA <= x"0010";
            when "10" & x"d32" => DATA <= x"0004";
            when "10" & x"d33" => DATA <= x"0028";
            when "10" & x"d34" => DATA <= x"e412";
            when "10" & x"d35" => DATA <= x"1904";
            when "10" & x"d36" => DATA <= x"f0cf";
            when "10" & x"d37" => DATA <= x"8000";
            when "10" & x"d38" => DATA <= x"2930";
            when "10" & x"d39" => DATA <= x"9a4c";
            when "10" & x"d3a" => DATA <= x"2252";
            when "10" & x"d3b" => DATA <= x"6137";
            when "10" & x"d3c" => DATA <= x"c03c";
            when "10" & x"d3d" => DATA <= x"03c0";
            when "10" & x"d3e" => DATA <= x"3800";
            when "10" & x"d3f" => DATA <= x"1140";
            when "10" & x"d40" => DATA <= x"008e";
            when "10" & x"d41" => DATA <= x"0004";
            when "10" & x"d42" => DATA <= x"7804";
            when "10" & x"d43" => DATA <= x"8008";
            when "10" & x"d44" => DATA <= x"3c03";
            when "10" & x"d45" => DATA <= x"4008";
            when "10" & x"d46" => DATA <= x"1400";
            when "10" & x"d47" => DATA <= x"40f0";
            when "10" & x"d48" => DATA <= x"0f00";
            when "10" & x"d49" => DATA <= x"f00f";
            when "10" & x"d4a" => DATA <= x"00f0";
            when "10" & x"d4b" => DATA <= x"0000";
            when "10" & x"d4c" => DATA <= x"0a80";
            when "10" & x"d4d" => DATA <= x"0040";
            when "10" & x"d4e" => DATA <= x"0017";
            when "10" & x"d4f" => DATA <= x"8078";
            when "10" & x"d50" => DATA <= x"0780";
            when "10" & x"d51" => DATA <= x"6800";
            when "10" & x"d52" => DATA <= x"4280";
            when "10" & x"d53" => DATA <= x"021e";
            when "10" & x"d54" => DATA <= x"01e0";
            when "10" & x"d55" => DATA <= x"1e01";
            when "10" & x"d56" => DATA <= x"e01f";
            when "10" & x"d57" => DATA <= x"0080";
            when "10" & x"d58" => DATA <= x"7e9f";
            when "10" & x"d59" => DATA <= x"5a8d";
            when "10" & x"d5a" => DATA <= x"d2a1";
            when "10" & x"d5b" => DATA <= x"70f8";
            when "10" & x"d5c" => DATA <= x"dc20";
            when "10" & x"d5d" => DATA <= x"5002";
            when "10" & x"d5e" => DATA <= x"cbc0";
            when "10" & x"d5f" => DATA <= x"2c00";
            when "10" & x"d60" => DATA <= x"a1c0";
            when "10" & x"d61" => DATA <= x"14a0";
            when "10" & x"d62" => DATA <= x"007f";
            when "10" & x"d63" => DATA <= x"8178";
            when "10" & x"d64" => DATA <= x"0003";
            when "10" & x"d65" => DATA <= x"4007";
            when "10" & x"d66" => DATA <= x"f057";
            when "10" & x"d67" => DATA <= x"0002";
            when "10" & x"d68" => DATA <= x"2802";
            when "10" & x"d69" => DATA <= x"8311";
            when "10" & x"d6a" => DATA <= x"9419";
            when "10" & x"d6b" => DATA <= x"c580";
            when "10" & x"d6c" => DATA <= x"0380";
            when "10" & x"d6d" => DATA <= x"1ce0";
            when "10" & x"d6e" => DATA <= x"0020";
            when "10" & x"d6f" => DATA <= x"153c";
            when "10" & x"d70" => DATA <= x"0380";
            when "10" & x"d71" => DATA <= x"040a";
            when "10" & x"d72" => DATA <= x"a100";
            when "10" & x"d73" => DATA <= x"0010";
            when "10" & x"d74" => DATA <= x"0010";
            when "10" & x"d75" => DATA <= x"0008";
            when "10" & x"d76" => DATA <= x"1c00";
            when "10" & x"d77" => DATA <= x"02e0";
            when "10" & x"d78" => DATA <= x"0200";
            when "10" & x"d79" => DATA <= x"5403";
            when "10" & x"d7a" => DATA <= x"c000";
            when "10" & x"d7b" => DATA <= x"4a0c";
            when "10" & x"d7c" => DATA <= x"0703";
            when "10" & x"d7d" => DATA <= x"0080";
            when "10" & x"d7e" => DATA <= x"ca04";
            when "10" & x"d7f" => DATA <= x"0020";
            when "10" & x"d80" => DATA <= x"2c00";
            when "10" & x"d81" => DATA <= x"0203";
            when "10" & x"d82" => DATA <= x"a010";
            when "10" & x"d83" => DATA <= x"0700";
            when "10" & x"d84" => DATA <= x"d085";
            when "10" & x"d85" => DATA <= x"0010";
            when "10" & x"d86" => DATA <= x"6400";
            when "10" & x"d87" => DATA <= x"03e0";
            when "10" & x"d88" => DATA <= x"028f";
            when "10" & x"d89" => DATA <= x"0060";
            when "10" & x"d8a" => DATA <= x"5803";
            when "10" & x"d8b" => DATA <= x"bd8e";
            when "10" & x"d8c" => DATA <= x"cf77";
            when "10" & x"d8d" => DATA <= x"f67a";
            when "10" & x"d8e" => DATA <= x"9d46";
            when "10" & x"d8f" => DATA <= x"ab54";
            when "10" & x"d90" => DATA <= x"a26a";
            when "10" & x"d91" => DATA <= x"8556";
            when "10" & x"d92" => DATA <= x"893f";
            when "10" & x"d93" => DATA <= x"9df9";
            when "10" & x"d94" => DATA <= x"fcbe";
            when "10" & x"d95" => DATA <= x"7f27";
            when "10" & x"d96" => DATA <= x"d608";
            when "10" & x"d97" => DATA <= x"e018";
            when "10" & x"d98" => DATA <= x"f800";
            when "10" & x"d99" => DATA <= x"0400";
            when "10" & x"d9a" => DATA <= x"03f0";
            when "10" & x"d9b" => DATA <= x"0a01";
            when "10" & x"d9c" => DATA <= x"f857";
            when "10" & x"d9d" => DATA <= x"9004";
            when "10" & x"d9e" => DATA <= x"277f";
            when "10" & x"d9f" => DATA <= x"b800";
            when "10" & x"da0" => DATA <= x"0c00";
            when "10" & x"da1" => DATA <= x"07ff";
            when "10" & x"da2" => DATA <= x"bfbf";
            when "10" & x"da3" => DATA <= x"fc03";
            when "10" & x"da4" => DATA <= x"6e21";
            when "10" & x"da5" => DATA <= x"10f0";
            when "10" & x"da6" => DATA <= x"72cd";
            when "10" & x"da7" => DATA <= x"3ffd";
            when "10" & x"da8" => DATA <= x"ff57";
            when "10" & x"da9" => DATA <= x"fc7e";
            when "10" & x"daa" => DATA <= x"0fa3";
            when "10" & x"dab" => DATA <= x"faff";
            when "10" & x"dac" => DATA <= x"afc9";
            when "10" & x"dad" => DATA <= x"003f";
            when "10" & x"dae" => DATA <= x"f7fc";
            when "10" & x"daf" => DATA <= x"8030";
            when "10" & x"db0" => DATA <= x"2b9d";
            when "10" & x"db1" => DATA <= x"9ee6";
            when "10" & x"db2" => DATA <= x"0057";
            when "10" & x"db3" => DATA <= x"005d";
            when "10" & x"db4" => DATA <= x"3e1b";
            when "10" & x"db5" => DATA <= x"0fa7";
            when "10" & x"db6" => DATA <= x"c3f5";
            when "10" & x"db7" => DATA <= x"3ed4";
            when "10" & x"db8" => DATA <= x"6ab5";
            when "10" & x"db9" => DATA <= x"198c";
            when "10" & x"dba" => DATA <= x"a64a";
            when "10" & x"dbb" => DATA <= x"2593";
            when "10" & x"dbc" => DATA <= x"feaf";
            when "10" & x"dbd" => DATA <= x"5f00";
            when "10" & x"dbe" => DATA <= x"f00a";
            when "10" & x"dbf" => DATA <= x"0002";
            when "10" & x"dc0" => DATA <= x"5000";
            when "10" & x"dc1" => DATA <= x"1280";
            when "10" & x"dc2" => DATA <= x"009e";
            when "10" & x"dc3" => DATA <= x"01e0";
            when "10" & x"dc4" => DATA <= x"1e01";
            when "10" & x"dc5" => DATA <= x"2002";
            when "10" & x"dc6" => DATA <= x"0a00";
            when "10" & x"dc7" => DATA <= x"1050";
            when "10" & x"dc8" => DATA <= x"0083";
            when "10" & x"dc9" => DATA <= x"c03c";
            when "10" & x"dca" => DATA <= x"03c0";
            when "10" & x"dcb" => DATA <= x"3c03";
            when "10" & x"dcc" => DATA <= x"c000";
            when "10" & x"dcd" => DATA <= x"001f";
            when "10" & x"dce" => DATA <= x"00f0";
            when "10" & x"dcf" => DATA <= x"0900";
            when "10" & x"dd0" => DATA <= x"0178";
            when "10" & x"dd1" => DATA <= x"0780";
            when "10" & x"dd2" => DATA <= x"0001";
            when "10" & x"dd3" => DATA <= x"1e01";
            when "10" & x"dd4" => DATA <= x"a001";
            when "10" & x"dd5" => DATA <= x"0a00";
            when "10" & x"dd6" => DATA <= x"0878";
            when "10" & x"dd7" => DATA <= x"0000";
            when "10" & x"dd8" => DATA <= x"1143";
            when "10" & x"dd9" => DATA <= x"209e";
            when "10" & x"dda" => DATA <= x"194c";
            when "10" & x"ddb" => DATA <= x"867c";
            when "10" & x"ddc" => DATA <= x"0001";
            when "10" & x"ddd" => DATA <= x"4984";
            when "10" & x"dde" => DATA <= x"4261";
            when "10" & x"ddf" => DATA <= x"108a";
            when "10" & x"de0" => DATA <= x"4c22";
            when "10" & x"de1" => DATA <= x"7807";
            when "10" & x"de2" => DATA <= x"8001";
            when "10" & x"de3" => DATA <= x"3c02";
            when "10" & x"de4" => DATA <= x"8001";
            when "10" & x"de5" => DATA <= x"1a00";
            when "10" & x"de6" => DATA <= x"08f0";
            when "10" & x"de7" => DATA <= x"0d00";
            when "10" & x"de8" => DATA <= x"1078";
            when "10" & x"de9" => DATA <= x"0780";
            when "10" & x"dea" => DATA <= x"0008";
            when "10" & x"deb" => DATA <= x"1e01";
            when "10" & x"dec" => DATA <= x"e01e";
            when "10" & x"ded" => DATA <= x"01e0";
            when "10" & x"dee" => DATA <= x"1e00";
            when "10" & x"def" => DATA <= x"0001";
            when "10" & x"df0" => DATA <= x"5000";
            when "10" & x"df1" => DATA <= x"0a80";
            when "10" & x"df2" => DATA <= x"005e";
            when "10" & x"df3" => DATA <= x"01e0";
            when "10" & x"df4" => DATA <= x"1e01";
            when "10" & x"df5" => DATA <= x"2001";
            when "10" & x"df6" => DATA <= x"0a00";
            when "10" & x"df7" => DATA <= x"0850";
            when "10" & x"df8" => DATA <= x"0043";
            when "10" & x"df9" => DATA <= x"c03c";
            when "10" & x"dfa" => DATA <= x"03c0";
            when "10" & x"dfb" => DATA <= x"2403";
            when "10" & x"dfc" => DATA <= x"e010";
            when "10" & x"dfd" => DATA <= x"0dc7";
            when "10" & x"dfe" => DATA <= x"e371";
            when "10" & x"dff" => DATA <= x"f81c";
            when "10" & x"e00" => DATA <= x"7a3f";
            when "10" & x"e01" => DATA <= x"1b80";
            when "10" & x"e02" => DATA <= x"0010";
            when "10" & x"e03" => DATA <= x"0004";
            when "10" & x"e04" => DATA <= x"6000";
            when "10" & x"e05" => DATA <= x"5207";
            when "10" & x"e06" => DATA <= x"8050";
            when "10" & x"e07" => DATA <= x"0050";
            when "10" & x"e08" => DATA <= x"8800";
            when "10" & x"e09" => DATA <= x"2800";
            when "10" & x"e0a" => DATA <= x"0a94";
            when "10" & x"e0b" => DATA <= x"0140";
            when "10" & x"e0c" => DATA <= x"200e";
            when "10" & x"e0d" => DATA <= x"01a0";
            when "10" & x"e0e" => DATA <= x"0100";
            when "10" & x"e0f" => DATA <= x"a000";
            when "10" & x"e10" => DATA <= x"0800";
            when "10" & x"e11" => DATA <= x"0880";
            when "10" & x"e12" => DATA <= x"02c0";
            when "10" & x"e13" => DATA <= x"40b1";
            when "10" & x"e14" => DATA <= x"580c";
            when "10" & x"e15" => DATA <= x"1603";
            when "10" & x"e16" => DATA <= x"0581";
            when "10" & x"e17" => DATA <= x"0a30";
            when "10" & x"e18" => DATA <= x"210c";
            when "10" & x"e19" => DATA <= x"2800";
            when "10" & x"e1a" => DATA <= x"0da0";
            when "10" & x"e1b" => DATA <= x"080e";
            when "10" & x"e1c" => DATA <= x"0051";
            when "10" & x"e1d" => DATA <= x"0204";
            when "10" & x"e1e" => DATA <= x"0000";
            when "10" & x"e1f" => DATA <= x"4000";
            when "10" & x"e20" => DATA <= x"41a0";
            when "10" & x"e21" => DATA <= x"040e";
            when "10" & x"e22" => DATA <= x"0028";
            when "10" & x"e23" => DATA <= x"0000";
            when "10" & x"e24" => DATA <= x"801e";
            when "10" & x"e25" => DATA <= x"00e0";
            when "10" & x"e26" => DATA <= x"c070";
            when "10" & x"e27" => DATA <= x"1283";
            when "10" & x"e28" => DATA <= x"00de";
            when "10" & x"e29" => DATA <= x"0000";
            when "10" & x"e2a" => DATA <= x"0480";
            when "10" & x"e2b" => DATA <= x"4060";
            when "10" & x"e2c" => DATA <= x"1007";
            when "10" & x"e2d" => DATA <= x"0095";
            when "10" & x"e2e" => DATA <= x"4005";
            when "10" & x"e2f" => DATA <= x"0020";
            when "10" & x"e30" => DATA <= x"0780";
            when "10" & x"e31" => DATA <= x"1400";
            when "10" & x"e32" => DATA <= x"0408";
            when "10" & x"e33" => DATA <= x"0003";
            when "10" & x"e34" => DATA <= x"4000";
            when "10" & x"e35" => DATA <= x"1050";
            when "10" & x"e36" => DATA <= x"0054";
            when "10" & x"e37" => DATA <= x"0041";
            when "10" & x"e38" => DATA <= x"5002";
            when "10" & x"e39" => DATA <= x"8000";
            when "10" & x"e3a" => DATA <= x"8060";
            when "10" & x"e3b" => DATA <= x"7002";
            when "10" & x"e3c" => DATA <= x"0001";
            when "10" & x"e3d" => DATA <= x"5cee";
            when "10" & x"e3e" => DATA <= x"36bb";
            when "10" & x"e3f" => DATA <= x"8d8e";
            when "10" & x"e40" => DATA <= x"e363";
            when "10" & x"e41" => DATA <= x"a2d0";
            when "10" & x"e42" => DATA <= x"0aa5";
            when "10" & x"e43" => DATA <= x"132b";
            when "10" & x"e44" => DATA <= x"aa9f";
            when "10" & x"e45" => DATA <= x"e7f3";
            when "10" & x"e46" => DATA <= x"dbfe";
            when "10" & x"e47" => DATA <= x"9fce";
            when "10" & x"e48" => DATA <= x"e7e7";
            when "10" & x"e49" => DATA <= x"0001";
            when "10" & x"e4a" => DATA <= x"1002";
            when "10" & x"e4b" => DATA <= x"7e3e";
            when "10" & x"e4c" => DATA <= x"0000";
            when "10" & x"e4d" => DATA <= x"102f";
            when "10" & x"e4e" => DATA <= x"003f";
            when "10" & x"e4f" => DATA <= x"c060";
            when "10" & x"e50" => DATA <= x"0705";
            when "10" & x"e51" => DATA <= x"4038";
            when "10" & x"e52" => DATA <= x"0c00";
            when "10" & x"e53" => DATA <= x"3002";
            when "10" & x"e54" => DATA <= x"391f";
            when "10" & x"e55" => DATA <= x"dfe0";
            when "10" & x"e56" => DATA <= x"1a00";
            when "10" & x"e57" => DATA <= x"9ff0";
            when "10" & x"e58" => DATA <= x"5b80";
            when "10" & x"e59" => DATA <= x"01df";
            when "10" & x"e5a" => DATA <= x"f402";
            when "10" & x"e5b" => DATA <= x"0000";
            when "10" & x"e5c" => DATA <= x"8038";
            when "10" & x"e5d" => DATA <= x"068d";
            when "10" & x"e5e" => DATA <= x"0614";
            when "10" & x"e5f" => DATA <= x"01c6";
            when "10" & x"e60" => DATA <= x"9dfe";
            when "10" & x"e61" => DATA <= x"0060";
            when "10" & x"e62" => DATA <= x"77ff";
            when "10" & x"e63" => DATA <= x"1f80";
            when "10" & x"e64" => DATA <= x"07fd";
            when "10" & x"e65" => DATA <= x"7f40";
            when "10" & x"e66" => DATA <= x"0fca";
            when "10" & x"e67" => DATA <= x"001f";
            when "10" & x"e68" => DATA <= x"bff8";
            when "10" & x"e69" => DATA <= x"02bf";
            when "10" & x"e6a" => DATA <= x"dc00";
            when "10" & x"e6b" => DATA <= x"07f8";
            when "10" & x"e6c" => DATA <= x"0080";
            when "10" & x"e6d" => DATA <= x"e667";
            when "10" & x"e6e" => DATA <= x"b1dc";
            when "10" & x"e6f" => DATA <= x"ec0a";
            when "10" & x"e70" => DATA <= x"e00f";
            when "10" & x"e71" => DATA <= x"a7c3";
            when "10" & x"e72" => DATA <= x"c1b4";
            when "10" & x"e73" => DATA <= x"f87c";
            when "10" & x"e74" => DATA <= x"3c1f";
            when "10" & x"e75" => DATA <= x"64b2";
            when "10" & x"e76" => DATA <= x"990c";
            when "10" & x"e77" => DATA <= x"062d";
            when "10" & x"e78" => DATA <= x"6230";
            when "10" & x"e79" => DATA <= x"27d5";
            when "10" & x"e7a" => DATA <= x"eef5";
            when "10" & x"e7b" => DATA <= x"af7b";
            when "10" & x"e7c" => DATA <= x"0022";
            when "10" & x"e7d" => DATA <= x"3cac";
            when "10" & x"e7e" => DATA <= x"0088";
            when "10" & x"e7f" => DATA <= x"f090";
            when "10" & x"e80" => DATA <= x"0e04";
            when "10" & x"e81" => DATA <= x"7078";
            when "10" & x"e82" => DATA <= x"0207";
            when "10" & x"e83" => DATA <= x"4028";
            when "10" & x"e84" => DATA <= x"2103";
            when "10" & x"e85" => DATA <= x"e008";
            when "10" & x"e86" => DATA <= x"6000";
            when "10" & x"e87" => DATA <= x"8280";
            when "10" & x"e88" => DATA <= x"3880";
            when "10" & x"e89" => DATA <= x"0760";
            when "10" & x"e8a" => DATA <= x"0400";
            when "10" & x"e8b" => DATA <= x"7e80";
            when "10" & x"e8c" => DATA <= x"5200";
            when "10" & x"e8d" => DATA <= x"3ec0";
            when "10" & x"e8e" => DATA <= x"0021";
            when "10" & x"e8f" => DATA <= x"cf00";
            when "10" & x"e90" => DATA <= x"0868";
            when "10" & x"e91" => DATA <= x"0500";
            when "10" & x"e92" => DATA <= x"9e2c";
            when "10" & x"e93" => DATA <= x"0044";
            when "10" & x"e94" => DATA <= x"78d0";
            when "10" & x"e95" => DATA <= x"0a02";
            when "10" & x"e96" => DATA <= x"7878";
            when "10" & x"e97" => DATA <= x"0383";
            when "10" & x"e98" => DATA <= x"4028";
            when "10" & x"e99" => DATA <= x"2181";
            when "10" & x"e9a" => DATA <= x"6000";
            when "10" & x"e9b" => DATA <= x"1018";
            when "10" & x"e9c" => DATA <= x"0021";
            when "10" & x"e9d" => DATA <= x"c001";
            when "10" & x"e9e" => DATA <= x"0088";
            when "10" & x"e9f" => DATA <= x"0f40";
            when "10" & x"ea0" => DATA <= x"1108";
            when "10" & x"ea1" => DATA <= x"e715";
            when "10" & x"ea2" => DATA <= x"0c82";
            when "10" & x"ea3" => DATA <= x"6865";
            when "10" & x"ea4" => DATA <= x"f8c0";
            when "10" & x"ea5" => DATA <= x"67e8";
            when "10" & x"ea6" => DATA <= x"03fc";
            when "10" & x"ea7" => DATA <= x"fe3f";
            when "10" & x"ea8" => DATA <= x"2693";
            when "10" & x"ea9" => DATA <= x"0884";
            when "10" & x"eaa" => DATA <= x"c26d";
            when "10" & x"eab" => DATA <= x"5f87";
            when "10" & x"eac" => DATA <= x"f400";
            when "10" & x"ead" => DATA <= x"0673";
            when "10" & x"eae" => DATA <= x"00e8";
            when "10" & x"eaf" => DATA <= x"0011";
            when "10" & x"eb0" => DATA <= x"0804";
            when "10" & x"eb1" => DATA <= x"b004";
            when "10" & x"eb2" => DATA <= x"4207";
            when "10" & x"eb3" => DATA <= x"4028";
            when "10" & x"eb4" => DATA <= x"2133";
            when "10" & x"eb5" => DATA <= x"e000";
            when "10" & x"eb6" => DATA <= x"3d00";
            when "10" & x"eb7" => DATA <= x"a201";
            when "10" & x"eb8" => DATA <= x"9580";
            when "10" & x"eb9" => DATA <= x"1001";
            when "10" & x"eba" => DATA <= x"a002";
            when "10" & x"ebb" => DATA <= x"0700";
            when "10" & x"ebc" => DATA <= x"7207";
            when "10" & x"ebd" => DATA <= x"8078";
            when "10" & x"ebe" => DATA <= x"0001";
            when "10" & x"ebf" => DATA <= x"21a0";
            when "10" & x"ec0" => DATA <= x"0011";
            when "10" & x"ec1" => DATA <= x"1966";
            when "10" & x"ec2" => DATA <= x"c004";
            when "10" & x"ec3" => DATA <= x"4600";
            when "10" & x"ec4" => DATA <= x"000a";
            when "10" & x"ec5" => DATA <= x"8038";
            when "10" & x"ec6" => DATA <= x"0905";
            when "10" & x"ec7" => DATA <= x"e008";
            when "10" & x"ec8" => DATA <= x"0d00";
            when "10" & x"ec9" => DATA <= x"0400";
            when "10" & x"eca" => DATA <= x"0196";
            when "10" & x"ecb" => DATA <= x"0011";
            when "10" & x"ecc" => DATA <= x"a000";
            when "10" & x"ecd" => DATA <= x"8500";
            when "10" & x"ece" => DATA <= x"5085";
            when "10" & x"ecf" => DATA <= x"08f8";
            when "10" & x"ed0" => DATA <= x"021f";
            when "10" & x"ed1" => DATA <= x"4004";
            when "10" & x"ed2" => DATA <= x"0aa3";
            when "10" & x"ed3" => DATA <= x"3580";
            when "10" & x"ed4" => DATA <= x"2000";
            when "10" & x"ed5" => DATA <= x"1b00";
            when "10" & x"ed6" => DATA <= x"40a8";
            when "10" & x"ed7" => DATA <= x"07e7";
            when "10" & x"ed8" => DATA <= x"6e07";
            when "10" & x"ed9" => DATA <= x"1bc9";
            when "10" & x"eda" => DATA <= x"e1f2";
            when "10" & x"edb" => DATA <= x"e000";
            when "10" & x"edc" => DATA <= x"0400";
            when "10" & x"edd" => DATA <= x"0d13";
            when "10" & x"ede" => DATA <= x"022a";
            when "10" & x"edf" => DATA <= x"00e8";
            when "10" & x"ee0" => DATA <= x"0601";
            when "10" & x"ee1" => DATA <= x"014b";
            when "10" & x"ee2" => DATA <= x"401c";
            when "10" & x"ee3" => DATA <= x"0200";
            when "10" & x"ee4" => DATA <= x"1494";
            when "10" & x"ee5" => DATA <= x"b800";
            when "10" & x"ee6" => DATA <= x"0340";
            when "10" & x"ee7" => DATA <= x"0016";
            when "10" & x"ee8" => DATA <= x"9700";
            when "10" & x"ee9" => DATA <= x"0838";
            when "10" & x"eea" => DATA <= x"0004";
            when "10" & x"eeb" => DATA <= x"8016";
            when "10" & x"eec" => DATA <= x"0338";
            when "10" & x"eed" => DATA <= x"b056";
            when "10" & x"eee" => DATA <= x"0804";
            when "10" & x"eef" => DATA <= x"8006";
            when "10" & x"ef0" => DATA <= x"0001";
            when "10" & x"ef1" => DATA <= x"8152";
            when "10" & x"ef2" => DATA <= x"8004";
            when "10" & x"ef3" => DATA <= x"1e00";
            when "10" & x"ef4" => DATA <= x"0045";
            when "10" & x"ef5" => DATA <= x"2200";
            when "10" & x"ef6" => DATA <= x"0a00";
            when "10" & x"ef7" => DATA <= x"0280";
            when "10" & x"ef8" => DATA <= x"008a";
            when "10" & x"ef9" => DATA <= x"f000";
            when "10" & x"efa" => DATA <= x"1004";
            when "10" & x"efb" => DATA <= x"2bc0";
            when "10" & x"efc" => DATA <= x"0050";
            when "10" & x"efd" => DATA <= x"0006";
            when "10" & x"efe" => DATA <= x"8300";
            when "10" & x"eff" => DATA <= x"80ca";
            when "10" & x"f00" => DATA <= x"04a0";
            when "10" & x"f01" => DATA <= x"cf00";
            when "10" & x"f02" => DATA <= x"4048";
            when "10" & x"f03" => DATA <= x"0802";
            when "10" & x"f04" => DATA <= x"8040";
            when "10" & x"f05" => DATA <= x"7200";
            when "10" & x"f06" => DATA <= x"0400";
            when "10" & x"f07" => DATA <= x"054a";
            when "10" & x"f08" => DATA <= x"9400";
            when "10" & x"f09" => DATA <= x"21e0";
            when "10" & x"f0a" => DATA <= x"0400";
            when "10" & x"f0b" => DATA <= x"0680";
            when "10" & x"f0c" => DATA <= x"0440";
            when "10" & x"f0d" => DATA <= x"0050";
            when "10" & x"f0e" => DATA <= x"0282";
            when "10" & x"f0f" => DATA <= x"b801";
            when "10" & x"f10" => DATA <= x"0140";
            when "10" & x"f11" => DATA <= x"0106";
            when "10" & x"f12" => DATA <= x"031d";
            when "10" & x"f13" => DATA <= x"86c7";
            when "10" & x"f14" => DATA <= x"61b1";
            when "10" & x"f15" => DATA <= x"daeb";
            when "10" & x"f16" => DATA <= x"f39a";
            when "10" & x"f17" => DATA <= x"0ba0";
            when "10" & x"f18" => DATA <= x"2a29";
            when "10" & x"f19" => DATA <= x"5080";
            when "10" & x"f1a" => DATA <= x"f7f2";
            when "10" & x"f1b" => DATA <= x"fb07";
            when "10" & x"f1c" => DATA <= x"c01f";
            when "10" & x"f1d" => DATA <= x"efce";
            when "10" & x"f1e" => DATA <= x"0002";
            when "10" & x"f1f" => DATA <= x"001f";
            when "10" & x"f20" => DATA <= x"88f4";
            when "10" & x"f21" => DATA <= x"1a00";
            when "10" & x"f22" => DATA <= x"0150";
            when "10" & x"f23" => DATA <= x"0004";
            when "10" & x"f24" => DATA <= x"2fff";
            when "10" & x"f25" => DATA <= x"fffd";
            when "10" & x"f26" => DATA <= x"7ff8";
            when "10" & x"f27" => DATA <= x"0807";
            when "10" & x"f28" => DATA <= x"4d28";
            when "10" & x"f29" => DATA <= x"d801";
            when "10" & x"f2a" => DATA <= x"7fe7";
            when "10" & x"f2b" => DATA <= x"f005";
            when "10" & x"f2c" => DATA <= x"5fd1";
            when "10" & x"f2d" => DATA <= x"fd5f";
            when "10" & x"f2e" => DATA <= x"f803";
            when "10" & x"f2f" => DATA <= x"ffc0";
            when "10" & x"f30" => DATA <= x"0fe7";
            when "10" & x"f31" => DATA <= x"8a00";
            when "10" & x"f32" => DATA <= x"ae26";
            when "10" & x"f33" => DATA <= x"1382";
            when "10" & x"f34" => DATA <= x"b01c";
            when "10" & x"f35" => DATA <= x"f43e";
            when "10" & x"f36" => DATA <= x"9fa1";
            when "10" & x"f37" => DATA <= x"f0f0";
            when "10" & x"f38" => DATA <= x"5d3e";
            when "10" & x"f39" => DATA <= x"01a8";
            when "10" & x"f3a" => DATA <= x"100a";
            when "10" & x"f3b" => DATA <= x"2068";
            when "10" & x"f3c" => DATA <= x"d06a";
            when "10" & x"f3d" => DATA <= x"bf1f";
            when "10" & x"f3e" => DATA <= x"afc7";
            when "10" & x"f3f" => DATA <= x"a4f8";
            when "10" & x"f40" => DATA <= x"0000";
            when "10" & x"f41" => DATA <= x"4001";
            when "10" & x"f42" => DATA <= x"e3f1";
            when "10" & x"f43" => DATA <= x"5600";
            when "10" & x"f44" => DATA <= x"0470";
            when "10" & x"f45" => DATA <= x"007d";
            when "10" & x"f46" => DATA <= x"feaf";
            when "10" & x"f47" => DATA <= x"a00a";
            when "10" & x"f48" => DATA <= x"0400";
            when "10" & x"f49" => DATA <= x"26df";
            when "10" & x"f4a" => DATA <= x"ebfd";
            when "10" & x"f4b" => DATA <= x"000e";
            when "10" & x"f4c" => DATA <= x"3fde";
            when "10" & x"f4d" => DATA <= x"7400";
            when "10" & x"f4e" => DATA <= x"100c";
            when "10" & x"f4f" => DATA <= x"0007";
            when "10" & x"f50" => DATA <= x"cff6";
            when "10" & x"f51" => DATA <= x"de80";
            when "10" & x"f52" => DATA <= x"0e1f";
            when "10" & x"f53" => DATA <= x"e6da";
            when "10" & x"f54" => DATA <= x"0010";
            when "10" & x"f55" => DATA <= x"0c00";
            when "10" & x"f56" => DATA <= x"0dda";
            when "10" & x"f57" => DATA <= x"ffd0";
            when "10" & x"f58" => DATA <= x"0723";
            when "10" & x"f59" => DATA <= x"fde3";
            when "10" & x"f5a" => DATA <= x"4004";
            when "10" & x"f5b" => DATA <= x"0600";
            when "10" & x"f5c" => DATA <= x"01e8";
            when "10" & x"f5d" => DATA <= x"ff78";
            when "10" & x"f5e" => DATA <= x"e803";
            when "10" & x"f5f" => DATA <= x"21fe";
            when "10" & x"f60" => DATA <= x"ead0";
            when "10" & x"f61" => DATA <= x"061b";
            when "10" & x"f62" => DATA <= x"fd77";
            when "10" & x"f63" => DATA <= x"4014";
            when "10" & x"f64" => DATA <= x"0200";
            when "10" & x"f65" => DATA <= x"433f";
            when "10" & x"f66" => DATA <= x"d9fa";
            when "10" & x"f67" => DATA <= x"0087";
            when "10" & x"f68" => DATA <= x"7fb3";
            when "10" & x"f69" => DATA <= x"e802";
            when "10" & x"f6a" => DATA <= x"8180";
            when "10" & x"f6b" => DATA <= x"04d7";
            when "10" & x"f6c" => DATA <= x"f97e";
            when "10" & x"f6d" => DATA <= x"80b8";
            when "10" & x"f6e" => DATA <= x"009c";
            when "10" & x"f6f" => DATA <= x"ff2f";
            when "10" & x"f70" => DATA <= x"d000";
            when "10" & x"f71" => DATA <= x"2018";
            when "10" & x"f72" => DATA <= x"0013";
            when "10" & x"f73" => DATA <= x"bfcf";
            when "10" & x"f74" => DATA <= x"fa00";
            when "10" & x"f75" => DATA <= x"1c7f";
            when "10" & x"f76" => DATA <= x"bba8";
            when "10" & x"f77" => DATA <= x"0284";
            when "10" & x"f78" => DATA <= x"000e";
            when "10" & x"f79" => DATA <= x"c7fb";
            when "10" & x"f7a" => DATA <= x"df80";
            when "10" & x"f7b" => DATA <= x"1814";
            when "10" & x"f7c" => DATA <= x"0002";
            when "10" & x"f7d" => DATA <= x"7fd0";
            when "10" & x"f7e" => DATA <= x"0031";
            when "10" & x"f7f" => DATA <= x"0208";
            when "10" & x"f80" => DATA <= x"1000";
            when "10" & x"f81" => DATA <= x"1ff4";
            when "10" & x"f82" => DATA <= x"0010";
            when "10" & x"f83" => DATA <= x"0388";
            when "10" & x"f84" => DATA <= x"2801";
            when "10" & x"f85" => DATA <= x"ffc0";
            when "10" & x"f86" => DATA <= x"07e7";
            when "10" & x"f87" => DATA <= x"0500";
            when "10" & x"f88" => DATA <= x"3fe8";
            when "10" & x"f89" => DATA <= x"0006";
            when "10" & x"f8a" => DATA <= x"e000";
            when "10" & x"f8b" => DATA <= x"5403";
            when "10" & x"f8c" => DATA <= x"fe98";
            when "10" & x"f8d" => DATA <= x"00c0";
            when "10" & x"f8e" => DATA <= x"7000";
            when "10" & x"f8f" => DATA <= x"6dfe";
            when "10" & x"f90" => DATA <= x"f7d0";
            when "10" & x"f91" => DATA <= x"02f3";
            when "10" & x"f92" => DATA <= x"fd37";
            when "10" & x"f93" => DATA <= x"4000";
            when "10" & x"f94" => DATA <= x"80c0";
            when "10" & x"f95" => DATA <= x"002c";
            when "10" & x"f96" => DATA <= x"ff6d";
            when "10" & x"f97" => DATA <= x"e800";
            when "10" & x"f98" => DATA <= x"e1fe";
            when "10" & x"f99" => DATA <= x"e5a0";
            when "10" & x"f9a" => DATA <= x"0100";
            when "10" & x"f9b" => DATA <= x"c000";
            when "10" & x"f9c" => DATA <= x"dd7f";
            when "10" & x"f9d" => DATA <= x"bf74";
            when "10" & x"f9e" => DATA <= x"01e6";
            when "10" & x"f9f" => DATA <= x"ff78";
            when "10" & x"fa0" => DATA <= x"f001";
            when "10" & x"fa1" => DATA <= x"0000";
            when "10" & x"fa2" => DATA <= x"b07f";
            when "10" & x"fa3" => DATA <= x"be34";
            when "10" & x"fa4" => DATA <= x"0190";
            when "10" & x"fa5" => DATA <= x"ff75";
            when "10" & x"fa6" => DATA <= x"f002";
            when "10" & x"fa7" => DATA <= x"0000";
            when "10" & x"fa8" => DATA <= x"c97f";
            when "10" & x"fa9" => DATA <= x"bae8";
            when "10" & x"faa" => DATA <= x"0280";
            when "10" & x"fab" => DATA <= x"400d";
            when "10" & x"fac" => DATA <= x"27fb";
            when "10" & x"fad" => DATA <= x"3f40";
            when "10" & x"fae" => DATA <= x"10ef";
            when "10" & x"faf" => DATA <= x"f6ed";
            when "10" & x"fb0" => DATA <= x"0050";
            when "10" & x"fb1" => DATA <= x"1000";
            when "10" & x"fb2" => DATA <= x"1aff";
            when "10" & x"fb3" => DATA <= x"3de8";
            when "10" & x"fb4" => DATA <= x"003d";
            when "10" & x"fb5" => DATA <= x"fe1f";
            when "10" & x"fb6" => DATA <= x"e000";
            when "10" & x"fb7" => DATA <= x"6000";
            when "10" & x"fb8" => DATA <= x"1cff";
            when "10" & x"fb9" => DATA <= x"5ee8";
            when "10" & x"fba" => DATA <= x"02f1";
            when "10" & x"fbb" => DATA <= x"feae";
            when "10" & x"fbc" => DATA <= x"a00a";
            when "10" & x"fbd" => DATA <= x"1000";
            when "10" & x"fbe" => DATA <= x"1b1f";
            when "10" & x"fbf" => DATA <= x"efe0";
            when "10" & x"fc0" => DATA <= x"00c3";
            when "10" & x"fc1" => DATA <= x"800e";
            when "10" & x"fc2" => DATA <= x"4ff7";
            when "10" & x"fc3" => DATA <= x"d800";
            when "10" & x"fc4" => DATA <= x"2620";
            when "10" & x"fc5" => DATA <= x"3000";
            when "10" & x"fc6" => DATA <= x"1e4f";
            when "10" & x"fc7" => DATA <= x"f7d6";
            when "10" & x"fc8" => DATA <= x"8039";
            when "10" & x"fc9" => DATA <= x"1fef";
            when "10" & x"fca" => DATA <= x"1d00";
            when "10" & x"fcb" => DATA <= x"203f";
            when "10" & x"fcc" => DATA <= x"d2a9";
            when "10" & x"fcd" => DATA <= x"8000";
            when "10" & x"fce" => DATA <= x"fa9f";
            when "10" & x"fcf" => DATA <= x"a9fc";
            when "10" & x"fd0" => DATA <= x"fcaf";
            when "10" & x"fd1" => DATA <= x"1f80";
            when "10" & x"fd2" => DATA <= x"41a4";
            when "10" & x"fd3" => DATA <= x"0070";
            when "10" & x"fd4" => DATA <= x"0120";
            when "10" & x"fd5" => DATA <= x"ff00";
            when "10" & x"fd6" => DATA <= x"809e";
            when "10" & x"fd7" => DATA <= x"e000";
            when "10" & x"fd8" => DATA <= x"1500";
            when "10" & x"fd9" => DATA <= x"3fe8";
            when "10" & x"fda" => DATA <= x"0033";
            when "10" & x"fdb" => DATA <= x"4000";
            when "10" & x"fdc" => DATA <= x"4203";
            when "10" & x"fdd" => DATA <= x"fc88";
            when "10" & x"fde" => DATA <= x"807f";
            when "10" & x"fdf" => DATA <= x"8198";
            when "10" & x"fe0" => DATA <= x"6f80";
            when "10" & x"fe1" => DATA <= x"03fc";
            when "10" & x"fe2" => DATA <= x"0080";
            when "10" & x"fe3" => DATA <= x"013b";
            when "10" & x"fe4" => DATA <= x"41e0";
            when "10" & x"fe5" => DATA <= x"300b";
            when "10" & x"fe6" => DATA <= x"fc00";
            when "10" & x"fe7" => DATA <= x"88a0";
            when "10" & x"fe8" => DATA <= x"f182";
            when "10" & x"fe9" => DATA <= x"d1e2";
            when "10" & x"fea" => DATA <= x"0f00";
            when "10" & x"feb" => DATA <= x"11c0";
            when "10" & x"fec" => DATA <= x"8000";
            when "10" & x"fed" => DATA <= x"8700";
            when "10" & x"fee" => DATA <= x"0228";
            when "10" & x"fef" => DATA <= x"06c0";
            when "10" & x"ff0" => DATA <= x"1542";
            when "10" & x"ff1" => DATA <= x"8d00";
            when "10" & x"ff2" => DATA <= x"1000";
            when "10" & x"ff3" => DATA <= x"0800";
            when "10" & x"ff4" => DATA <= x"000d";
            when "10" & x"ff5" => DATA <= x"0007";
            when "10" & x"ff6" => DATA <= x"8094";
            when "10" & x"ff7" => DATA <= x"2ba0";
            when "10" & x"ff8" => DATA <= x"0040";
            when "10" & x"ff9" => DATA <= x"7031";
            when "10" & x"ffa" => DATA <= x"f9e0";
            when "10" & x"ffb" => DATA <= x"0ffe";
            when "10" & x"ffc" => DATA <= x"00a8";
            when "10" & x"ffd" => DATA <= x"0a01";
            when "10" & x"ffe" => DATA <= x"02c8";
            when "10" & x"fff" => DATA <= x"000c";
            when "11" & x"000" => DATA <= x"a010";
            when "11" & x"001" => DATA <= x"4078";
            when "11" & x"002" => DATA <= x"000b";
            when "11" & x"003" => DATA <= x"8000";
            when "11" & x"004" => DATA <= x"4000";
            when "11" & x"005" => DATA <= x"5700";
            when "11" & x"006" => DATA <= x"2815";
            when "11" & x"007" => DATA <= x"5200";
            when "11" & x"008" => DATA <= x"a0ae";
            when "11" & x"009" => DATA <= x"a742";
            when "11" & x"00a" => DATA <= x"0000";
            when "11" & x"00b" => DATA <= x"f339";
            when "11" & x"00c" => DATA <= x"d799";
            when "11" & x"00d" => DATA <= x"cde6";
            when "11" & x"00e" => DATA <= x"6321";
            when "11" & x"00f" => DATA <= x"a094";
            when "11" & x"010" => DATA <= x"5d54";
            when "11" & x"011" => DATA <= x"8a44";
            when "11" & x"012" => DATA <= x"202d";
            when "11" & x"013" => DATA <= x"fc8e";
            when "11" & x"014" => DATA <= x"7f00";
            when "11" & x"015" => DATA <= x"3158";
            when "11" & x"016" => DATA <= x"2380";
            when "11" & x"017" => DATA <= x"c3e0";
            when "11" & x"018" => DATA <= x"0010";
            when "11" & x"019" => DATA <= x"7e3f";
            when "11" & x"01a" => DATA <= x"c060";
            when "11" & x"01b" => DATA <= x"0783";
            when "11" & x"01c" => DATA <= x"fe80";
            when "11" & x"01d" => DATA <= x"1020";
            when "11" & x"01e" => DATA <= x"7003";
            when "11" & x"01f" => DATA <= x"fabf";
            when "11" & x"020" => DATA <= x"dc08";
            when "11" & x"021" => DATA <= x"007b";
            when "11" & x"022" => DATA <= x"8001";
            when "11" & x"023" => DATA <= x"bfe8";
            when "11" & x"024" => DATA <= x"07fb";
            when "11" & x"025" => DATA <= x"437f";
            when "11" & x"026" => DATA <= x"ec06";
            when "11" & x"027" => DATA <= x"9040";
            when "11" & x"028" => DATA <= x"1468";
            when "11" & x"029" => DATA <= x"36a3";
            when "11" & x"02a" => DATA <= x"4a36";
            when "11" & x"02b" => DATA <= x"7a7f";
            when "11" & x"02c" => DATA <= x"ff1f";
            when "11" & x"02d" => DATA <= x"83e4";
            when "11" & x"02e" => DATA <= x"febf";
            when "11" & x"02f" => DATA <= x"3c01";
            when "11" & x"030" => DATA <= x"ff60";
            when "11" & x"031" => DATA <= x"0e66";
            when "11" & x"032" => DATA <= x"7b98";
            when "11" & x"033" => DATA <= x"015c";
            when "11" & x"034" => DATA <= x"0407";
            when "11" & x"035" => DATA <= x"706c";
            when "11" & x"036" => DATA <= x"3e9f";
            when "11" & x"037" => DATA <= x"0fd4";
            when "11" & x"038" => DATA <= x"f87d";
            when "11" & x"039" => DATA <= x"3ed5";
            when "11" & x"03a" => DATA <= x"6837";
            when "11" & x"03b" => DATA <= x"1baf";
            when "11" & x"03c" => DATA <= x"53eb";
            when "11" & x"03d" => DATA <= x"e4e0";
            when "11" & x"03e" => DATA <= x"f4ef";
            when "11" & x"03f" => DATA <= x"078b";
            when "11" & x"040" => DATA <= x"cebf";
            when "11" & x"041" => DATA <= x"d803";
            when "11" & x"042" => DATA <= x"0002";
            when "11" & x"043" => DATA <= x"0160";
            when "11" & x"044" => DATA <= x"340a";
            when "11" & x"045" => DATA <= x"031a";
            when "11" & x"046" => DATA <= x"c00a";
            when "11" & x"047" => DATA <= x"1049";
            when "11" & x"048" => DATA <= x"b416";
            when "11" & x"049" => DATA <= x"0e30";
            when "11" & x"04a" => DATA <= x"08d0";
            when "11" & x"04b" => DATA <= x"e844";
            when "11" & x"04c" => DATA <= x"002e";
            when "11" & x"04d" => DATA <= x"2bfe";
            when "11" & x"04e" => DATA <= x"8100";
            when "11" & x"04f" => DATA <= x"0fc0";
            when "11" & x"050" => DATA <= x"03de";
            when "11" & x"051" => DATA <= x"bff8";
            when "11" & x"052" => DATA <= x"01fc";
            when "11" & x"053" => DATA <= x"b87f";
            when "11" & x"054" => DATA <= x"aede";
            when "11" & x"055" => DATA <= x"5400";
            when "11" & x"056" => DATA <= x"8006";
            when "11" & x"057" => DATA <= x"9e88";
            when "11" & x"058" => DATA <= x"04a6";
            when "11" & x"059" => DATA <= x"5001";
            when "11" & x"05a" => DATA <= x"2efe";
            when "11" & x"05b" => DATA <= x"4438";
            when "11" & x"05c" => DATA <= x"7bbc";
            when "11" & x"05d" => DATA <= x"00b4";
            when "11" & x"05e" => DATA <= x"7abf";
            when "11" & x"05f" => DATA <= x"eaf4";
            when "11" & x"060" => DATA <= x"7e3d";
            when "11" & x"061" => DATA <= x"a002";
            when "11" & x"062" => DATA <= x"dd3d";
            when "11" & x"063" => DATA <= x"8280";
            when "11" & x"064" => DATA <= x"5c00";
            when "11" & x"065" => DATA <= x"07d0";
            when "11" & x"066" => DATA <= x"0aa0";
            when "11" & x"067" => DATA <= x"583e";
            when "11" & x"068" => DATA <= x"2400";
            when "11" & x"069" => DATA <= x"8280";
            when "11" & x"06a" => DATA <= x"1800";
            when "11" & x"06b" => DATA <= x"5a1c";
            when "11" & x"06c" => DATA <= x"0004";
            when "11" & x"06d" => DATA <= x"04b0";
            when "11" & x"06e" => DATA <= x"0000";
            when "11" & x"06f" => DATA <= x"a415";
            when "11" & x"070" => DATA <= x"0000";
            when "11" & x"071" => DATA <= x"814d";
            when "11" & x"072" => DATA <= x"0602";
            when "11" & x"073" => DATA <= x"8421";
            when "11" & x"074" => DATA <= x"c00d";
            when "11" & x"075" => DATA <= x"00bb";
            when "11" & x"076" => DATA <= x"0000";
            when "11" & x"077" => DATA <= x"04e0";
            when "11" & x"078" => DATA <= x"0398";
            when "11" & x"079" => DATA <= x"55c0";
            when "11" & x"07a" => DATA <= x"0390";
            when "11" & x"07b" => DATA <= x"0728";
            when "11" & x"07c" => DATA <= x"d454";
            when "11" & x"07d" => DATA <= x"fbe0";
            when "11" & x"07e" => DATA <= x"0300";
            when "11" & x"07f" => DATA <= x"e380";
            when "11" & x"080" => DATA <= x"7800";
            when "11" & x"081" => DATA <= x"1415";
            when "11" & x"082" => DATA <= x"e001";
            when "11" & x"083" => DATA <= x"4700";
            when "11" & x"084" => DATA <= x"0228";
            when "11" & x"085" => DATA <= x"0281";
            when "11" & x"086" => DATA <= x"2800";
            when "11" & x"087" => DATA <= x"1415";
            when "11" & x"088" => DATA <= x"e000";
            when "11" & x"089" => DATA <= x"2500";
            when "11" & x"08a" => DATA <= x"0a8a";
            when "11" & x"08b" => DATA <= x"b600";
            when "11" & x"08c" => DATA <= x"3c18";
            when "11" & x"08d" => DATA <= x"0a0c";
            when "11" & x"08e" => DATA <= x"0c27";
            when "11" & x"08f" => DATA <= x"d508";
            when "11" & x"090" => DATA <= x"7001";
            when "11" & x"091" => DATA <= x"5280";
            when "11" & x"092" => DATA <= x"6c00";
            when "11" & x"093" => DATA <= x"de0e";
            when "11" & x"094" => DATA <= x"2718";
            when "11" & x"095" => DATA <= x"3801";
            when "11" & x"096" => DATA <= x"fe03";
            when "11" & x"097" => DATA <= x"0080";
            when "11" & x"098" => DATA <= x"005c";
            when "11" & x"099" => DATA <= x"00ff";
            when "11" & x"09a" => DATA <= x"a04d";
            when "11" & x"09b" => DATA <= x"007f";
            when "11" & x"09c" => DATA <= x"e800";
            when "11" & x"09d" => DATA <= x"8004";
            when "11" & x"09e" => DATA <= x"ffb0";
            when "11" & x"09f" => DATA <= x"0183";
            when "11" & x"0a0" => DATA <= x"fe82";
            when "11" & x"0a1" => DATA <= x"3801";
            when "11" & x"0a2" => DATA <= x"800d";
            when "11" & x"0a3" => DATA <= x"7f88";
            when "11" & x"0a4" => DATA <= x"2401";
            when "11" & x"0a5" => DATA <= x"8e00";
            when "11" & x"0a6" => DATA <= x"7fe8";
            when "11" & x"0a7" => DATA <= x"000c";
            when "11" & x"0a8" => DATA <= x"84ff";
            when "11" & x"0a9" => DATA <= x"0091";
            when "11" & x"0aa" => DATA <= x"3800";
            when "11" & x"0ab" => DATA <= x"c000";
            when "11" & x"0ac" => DATA <= x"7ff0";
            when "11" & x"0ad" => DATA <= x"0008";
            when "11" & x"0ae" => DATA <= x"0003";
            when "11" & x"0af" => DATA <= x"003f";
            when "11" & x"0b0" => DATA <= x"e800";
            when "11" & x"0b1" => DATA <= x"0200";
            when "11" & x"0b2" => DATA <= x"0110";
            when "11" & x"0b3" => DATA <= x"900f";
            when "11" & x"0b4" => DATA <= x"fd00";
            when "11" & x"0b5" => DATA <= x"00b0";
            when "11" & x"0b6" => DATA <= x"5ff3";
            when "11" & x"0b7" => DATA <= x"c140";
            when "11" & x"0b8" => DATA <= x"0c9e";
            when "11" & x"0b9" => DATA <= x"cb25";
            when "11" & x"0ba" => DATA <= x"0228";
            when "11" & x"0bb" => DATA <= x"0004";
            when "11" & x"0bc" => DATA <= x"05a0";
            when "11" & x"0bd" => DATA <= x"1027";
            when "11" & x"0be" => DATA <= x"003c";
            when "11" & x"0bf" => DATA <= x"1815";
            when "11" & x"0c0" => DATA <= x"0010";
            when "11" & x"0c1" => DATA <= x"e00a";
            when "11" & x"0c2" => DATA <= x"0100";
            when "11" & x"0c3" => DATA <= x"560b";
            when "11" & x"0c4" => DATA <= x"0380";
            when "11" & x"0c5" => DATA <= x"2a03";
            when "11" & x"0c6" => DATA <= x"403a";
            when "11" & x"0c7" => DATA <= x"0180";
            when "11" & x"0c8" => DATA <= x"f07b";
            when "11" & x"0c9" => DATA <= x"af47";
            when "11" & x"0ca" => DATA <= x"c8f0";
            when "11" & x"0cb" => DATA <= x"1b7d";
            when "11" & x"0cc" => DATA <= x"a2e3";
            when "11" & x"0cd" => DATA <= x"3416";
            when "11" & x"0ce" => DATA <= x"432f";
            when "11" & x"0cf" => DATA <= x"900b";
            when "11" & x"0d0" => DATA <= x"f5e0";
            when "11" & x"0d1" => DATA <= x"f13f";
            when "11" & x"0d2" => DATA <= x"9bc5";
            when "11" & x"0d3" => DATA <= x"6efe";
            when "11" & x"0d4" => DATA <= x"f070";
            when "11" & x"0d5" => DATA <= x"3c01";
            when "11" & x"0d6" => DATA <= x"a100";
            when "11" & x"0d7" => DATA <= x"2702";
            when "11" & x"0d8" => DATA <= x"bd87";
            when "11" & x"0d9" => DATA <= x"f608";
            when "11" & x"0da" => DATA <= x"b400";
            when "11" & x"0db" => DATA <= x"0438";
            when "11" & x"0dc" => DATA <= x"0283";
            when "11" & x"0dd" => DATA <= x"0afa";
            when "11" & x"0de" => DATA <= x"0141";
            when "11" & x"0df" => DATA <= x"03b0";
            when "11" & x"0e0" => DATA <= x"1821";
            when "11" & x"0e1" => DATA <= x"71d5";
            when "11" & x"0e2" => DATA <= x"0081";
            when "11" & x"0e3" => DATA <= x"7830";
            when "11" & x"0e4" => DATA <= x"00f7";
            when "11" & x"0e5" => DATA <= x"6abd";
            when "11" & x"0e6" => DATA <= x"1fe0";
            when "11" & x"0e7" => DATA <= x"07a3";
            when "11" & x"0e8" => DATA <= x"e040";
            when "11" & x"0e9" => DATA <= x"2ba2";
            when "11" & x"0ea" => DATA <= x"f379";
            when "11" & x"0eb" => DATA <= x"009e";
            when "11" & x"0ec" => DATA <= x"7f60";
            when "11" & x"0ed" => DATA <= x"0025";
            when "11" & x"0ee" => DATA <= x"00b2";
            when "11" & x"0ef" => DATA <= x"5c20";
            when "11" & x"0f0" => DATA <= x"0448";
            when "11" & x"0f1" => DATA <= x"000a";
            when "11" & x"0f2" => DATA <= x"402c";
            when "11" & x"0f3" => DATA <= x"9600";
            when "11" & x"0f4" => DATA <= x"001a";
            when "11" & x"0f5" => DATA <= x"00a4";
            when "11" & x"0f6" => DATA <= x"07d8";
            when "11" & x"0f7" => DATA <= x"52e0";
            when "11" & x"0f8" => DATA <= x"164b";
            when "11" & x"0f9" => DATA <= x"1b01";
            when "11" & x"0fa" => DATA <= x"0180";
            when "11" & x"0fb" => DATA <= x"7800";
            when "11" & x"0fc" => DATA <= x"2140";
            when "11" & x"0fd" => DATA <= x"0552";
            when "11" & x"0fe" => DATA <= x"0580";
            when "11" & x"0ff" => DATA <= x"2850";
            when "11" & x"100" => DATA <= x"2001";
            when "11" & x"101" => DATA <= x"0000";
            when "11" & x"102" => DATA <= x"0400";
            when "11" & x"103" => DATA <= x"050a";
            when "11" & x"104" => DATA <= x"9456";
            when "11" & x"105" => DATA <= x"0040";
            when "11" & x"106" => DATA <= x"0030";
            when "11" & x"107" => DATA <= x"9048";
            when "11" & x"108" => DATA <= x"3015";
            when "11" & x"109" => DATA <= x"4122";
            when "11" & x"10a" => DATA <= x"d068";
            when "11" & x"10b" => DATA <= x"8457";
            when "11" & x"10c" => DATA <= x"4054";
            when "11" & x"10d" => DATA <= x"52a8";
            when "11" & x"10e" => DATA <= x"9f4f";
            when "11" & x"10f" => DATA <= x"e7b7";
            when "11" & x"110" => DATA <= x"fd3f";
            when "11" & x"111" => DATA <= x"95c0";
            when "11" & x"112" => DATA <= x"0f10";
            when "11" & x"113" => DATA <= x"0a20";
            when "11" & x"114" => DATA <= x"04fc";
            when "11" & x"115" => DATA <= x"7c50";
            when "11" & x"116" => DATA <= x"000c";
            when "11" & x"117" => DATA <= x"0001";
            when "11" & x"118" => DATA <= x"003f";
            when "11" & x"119" => DATA <= x"c1e0";
            when "11" & x"11a" => DATA <= x"0202";
            when "11" & x"11b" => DATA <= x"0000";
            when "11" & x"11c" => DATA <= x"e970";
            when "11" & x"11d" => DATA <= x"1fe8";
            when "11" & x"11e" => DATA <= x"037f";
            when "11" & x"11f" => DATA <= x"c066";
            when "11" & x"120" => DATA <= x"0006";
            when "11" & x"121" => DATA <= x"ffb8";
            when "11" & x"122" => DATA <= x"1fa5";
            when "11" & x"123" => DATA <= x"8009";
            when "11" & x"124" => DATA <= x"06c0";
            when "11" & x"125" => DATA <= x"4683";
            when "11" & x"126" => DATA <= x"6e00";
            when "11" & x"127" => DATA <= x"1851";
            when "11" & x"128" => DATA <= x"b57f";
            when "11" & x"129" => DATA <= x"d004";
            when "11" & x"12a" => DATA <= x"ff8f";
            when "11" & x"12b" => DATA <= x"c020";
            when "11" & x"12c" => DATA <= x"05f4";
            when "11" & x"12d" => DATA <= x"dfbf";
            when "11" & x"12e" => DATA <= x"2802";
            when "11" & x"12f" => DATA <= x"bff8";
            when "11" & x"130" => DATA <= x"01fe";
            when "11" & x"131" => DATA <= x"fc40";
            when "11" & x"132" => DATA <= x"001f";
            when "11" & x"133" => DATA <= x"fc00";
            when "11" & x"134" => DATA <= x"cf63";
            when "11" & x"135" => DATA <= x"b9d8";
            when "11" & x"136" => DATA <= x"15c0";
            when "11" & x"137" => DATA <= x"0070";
            when "11" & x"138" => DATA <= x"07c3";
            when "11" & x"139" => DATA <= x"69f0";
            when "11" & x"13a" => DATA <= x"f878";
            when "11" & x"13b" => DATA <= x"3e1e";
            when "11" & x"13c" => DATA <= x"0f86";
            when "11" & x"13d" => DATA <= x"0a80";
            when "11" & x"13e" => DATA <= x"5a46";
            when "11" & x"13f" => DATA <= x"2456";
            when "11" & x"140" => DATA <= x"2be5";
            when "11" & x"141" => DATA <= x"fee0";
            when "11" & x"142" => DATA <= x"0400";
            when "11" & x"143" => DATA <= x"1ff5";
            when "11" & x"144" => DATA <= x"7e01";
            when "11" & x"145" => DATA <= x"659f";
            when "11" & x"146" => DATA <= x"cf07";
            when "11" & x"147" => DATA <= x"07e3";
            when "11" & x"148" => DATA <= x"ddec";
            when "11" & x"149" => DATA <= x"4c7f";
            when "11" & x"14a" => DATA <= x"d803";
            when "11" & x"14b" => DATA <= x"89fd";
            when "11" & x"14c" => DATA <= x"200e";
            when "11" & x"14d" => DATA <= x"0783";
            when "11" & x"14e" => DATA <= x"5ddf";
            when "11" & x"14f" => DATA <= x"c00e";
            when "11" & x"150" => DATA <= x"a351";
            when "11" & x"151" => DATA <= x"2ea1";
            when "11" & x"152" => DATA <= x"b808";
            when "11" & x"153" => DATA <= x"0cfe";
            when "11" & x"154" => DATA <= x"6552";
            when "11" & x"155" => DATA <= x"5c80";
            when "11" & x"156" => DATA <= x"0040";
            when "11" & x"157" => DATA <= x"15df";
            when "11" & x"158" => DATA <= x"21c0";
            when "11" & x"159" => DATA <= x"3005";
            when "11" & x"15a" => DATA <= x"1ed8";
            when "11" & x"15b" => DATA <= x"0032";
            when "11" & x"15c" => DATA <= x"4010";
            when "11" & x"15d" => DATA <= x"0f00";
            when "11" & x"15e" => DATA <= x"2700";
            when "11" & x"15f" => DATA <= x"3004";
            when "11" & x"160" => DATA <= x"0007";
            when "11" & x"161" => DATA <= x"79e8";
            when "11" & x"162" => DATA <= x"403c";
            when "11" & x"163" => DATA <= x"000e";
            when "11" & x"164" => DATA <= x"47e0";
            when "11" & x"165" => DATA <= x"07fb";
            when "11" & x"166" => DATA <= x"0780";
            when "11" & x"167" => DATA <= x"1014";
            when "11" & x"168" => DATA <= x"0080";
            when "11" & x"169" => DATA <= x"0020";
            when "11" & x"16a" => DATA <= x"2801";
            when "11" & x"16b" => DATA <= x"0140";
            when "11" & x"16c" => DATA <= x"0800";
            when "11" & x"16d" => DATA <= x"0143";
            when "11" & x"16e" => DATA <= x"c028";
            when "11" & x"16f" => DATA <= x"0009";
            when "11" & x"170" => DATA <= x"a000";
            when "11" & x"171" => DATA <= x"8f00";
            when "11" & x"172" => DATA <= x"f00f";
            when "11" & x"173" => DATA <= x"00f0";
            when "11" & x"174" => DATA <= x"0e00";
            when "11" & x"175" => DATA <= x"2250";
            when "11" & x"176" => DATA <= x"0012";
            when "11" & x"177" => DATA <= x"8000";
            when "11" & x"178" => DATA <= x"8000";
            when "11" & x"179" => DATA <= x"2780";
            when "11" & x"17a" => DATA <= x"017c";
            when "11" & x"17b" => DATA <= x"0030";
            when "11" & x"17c" => DATA <= x"1048";
            when "11" & x"17d" => DATA <= x"0628";
            when "11" & x"17e" => DATA <= x"4030";
            when "11" & x"17f" => DATA <= x"10a0";
            when "11" & x"180" => DATA <= x"0058";
            when "11" & x"181" => DATA <= x"0a80";
            when "11" & x"182" => DATA <= x"0600";
            when "11" & x"183" => DATA <= x"0140";
            when "11" & x"184" => DATA <= x"0002";
            when "11" & x"185" => DATA <= x"13f0";
            when "11" & x"186" => DATA <= x"0d00";
            when "11" & x"187" => DATA <= x"0250";
            when "11" & x"188" => DATA <= x"0012";
            when "11" & x"189" => DATA <= x"8000";
            when "11" & x"18a" => DATA <= x"9e01";
            when "11" & x"18b" => DATA <= x"4002";
            when "11" & x"18c" => DATA <= x"0f00";
            when "11" & x"18d" => DATA <= x"e000";
            when "11" & x"18e" => DATA <= x"4500";
            when "11" & x"18f" => DATA <= x"023c";
            when "11" & x"190" => DATA <= x"0041";
            when "11" & x"191" => DATA <= x"e014";
            when "11" & x"192" => DATA <= x"0095";
            when "11" & x"193" => DATA <= x"0004";
            when "11" & x"194" => DATA <= x"0234";
            when "11" & x"195" => DATA <= x"0001";
            when "11" & x"196" => DATA <= x"f00e";
            when "11" & x"197" => DATA <= x"0010";
            when "11" & x"198" => DATA <= x"807c";
            when "11" & x"199" => DATA <= x"0340";
            when "11" & x"19a" => DATA <= x"021d";
            when "11" & x"19b" => DATA <= x"c000";
            when "11" & x"19c" => DATA <= x"1050";
            when "11" & x"19d" => DATA <= x"0081";
            when "11" & x"19e" => DATA <= x"f8fd";
            when "11" & x"19f" => DATA <= x"7f80";
            when "11" & x"1a0" => DATA <= x"0214";
            when "11" & x"1a1" => DATA <= x"0010";
            when "11" & x"1a2" => DATA <= x"4fd7";
            when "11" & x"1a3" => DATA <= x"fe80";
            when "11" & x"1a4" => DATA <= x"3993";
            when "11" & x"1a5" => DATA <= x"eff0";
            when "11" & x"1a6" => DATA <= x"0013";
            when "11" & x"1a7" => DATA <= x"803b";
            when "11" & x"1a8" => DATA <= x"fc00";
            when "11" & x"1a9" => DATA <= x"20a0";
            when "11" & x"1aa" => DATA <= x"0100";
            when "11" & x"1ab" => DATA <= x"02bf";
            when "11" & x"1ac" => DATA <= x"f401";
            when "11" & x"1ad" => DATA <= x"cebf";
            when "11" & x"1ae" => DATA <= x"7fc8";
            when "11" & x"1af" => DATA <= x"0009";
            when "11" & x"1b0" => DATA <= x"da9f";
            when "11" & x"1b1" => DATA <= x"7fe8";
            when "11" & x"1b2" => DATA <= x"010d";
            when "11" & x"1b3" => DATA <= x"067f";
            when "11" & x"1b4" => DATA <= x"d60a";
            when "11" & x"1b5" => DATA <= x"007a";
            when "11" & x"1b6" => DATA <= x"f802";
            when "11" & x"1b7" => DATA <= x"f740";
            when "11" & x"1b8" => DATA <= x"0040";
            when "11" & x"1b9" => DATA <= x"001f";
            when "11" & x"1ba" => DATA <= x"8058";
            when "11" & x"1bb" => DATA <= x"00f0";
            when "11" & x"1bc" => DATA <= x"005f";
            when "11" & x"1bd" => DATA <= x"d000";
            when "11" & x"1be" => DATA <= x"63b0";
            when "11" & x"1bf" => DATA <= x"1741";
            when "11" & x"1c0" => DATA <= x"0f8a";
            when "11" & x"1c1" => DATA <= x"007e";
            when "11" & x"1c2" => DATA <= x"bff8";
            when "11" & x"1c3" => DATA <= x"01fe";
            when "11" & x"1c4" => DATA <= x"0040";
            when "11" & x"1c5" => DATA <= x"1fcb";
            when "11" & x"1c6" => DATA <= x"fc00";
            when "11" & x"1c7" => DATA <= x"ff00";
            when "11" & x"1c8" => DATA <= x"0fc3";
            when "11" & x"1c9" => DATA <= x"8783";
            when "11" & x"1ca" => DATA <= x"e500";
            when "11" & x"1cb" => DATA <= x"3fc0";
            when "11" & x"1cc" => DATA <= x"0f46";
            when "11" & x"1cd" => DATA <= x"c0a2";
            when "11" & x"1ce" => DATA <= x"be00";
            when "11" & x"1cf" => DATA <= x"03f1";
            when "11" & x"1d0" => DATA <= x"c1e5";
            when "11" & x"1d1" => DATA <= x"e8b0";
            when "11" & x"1d2" => DATA <= x"5a3d";
            when "11" & x"1d3" => DATA <= x"1e14";
            when "11" & x"1d4" => DATA <= x"008e";
            when "11" & x"1d5" => DATA <= x"48a0";
            when "11" & x"1d6" => DATA <= x"5e07";
            when "11" & x"1d7" => DATA <= x"1700";
            when "11" & x"1d8" => DATA <= x"c280";
            when "11" & x"1d9" => DATA <= x"002f";
            when "11" & x"1da" => DATA <= x"f008";
            when "11" & x"1db" => DATA <= x"0006";
            when "11" & x"1dc" => DATA <= x"0200";
            when "11" & x"1dd" => DATA <= x"0880";
            when "11" & x"1de" => DATA <= x"0ffa";
            when "11" & x"1df" => DATA <= x"0070";
            when "11" & x"1e0" => DATA <= x"3e38";
            when "11" & x"1e1" => DATA <= x"01ff";
            when "11" & x"1e2" => DATA <= x"4014";
            when "11" & x"1e3" => DATA <= x"fe00";
            when "11" & x"1e4" => DATA <= x"7a00";
            when "11" & x"1e5" => DATA <= x"1ff4";
            when "11" & x"1e6" => DATA <= x"0040";
            when "11" & x"1e7" => DATA <= x"0052";
            when "11" & x"1e8" => DATA <= x"0001";
            when "11" & x"1e9" => DATA <= x"ff50";
            when "11" & x"1ea" => DATA <= x"0143";
            when "11" & x"1eb" => DATA <= x"2210";
            when "11" & x"1ec" => DATA <= x"a80a";
            when "11" & x"1ed" => DATA <= x"47b4";
            when "11" & x"1ee" => DATA <= x"5128";
            when "11" & x"1ef" => DATA <= x"8402";
            when "11" & x"1f0" => DATA <= x"2582";
            when "11" & x"1f1" => DATA <= x"aa41";
            when "11" & x"1f2" => DATA <= x"206a";
            when "11" & x"1f3" => DATA <= x"aaa0";
            when "11" & x"1f4" => DATA <= x"9567";
            when "11" & x"1f5" => DATA <= x"ef7f";
            when "11" & x"1f6" => DATA <= x"00b1";
            when "11" & x"1f7" => DATA <= x"6800";
            when "11" & x"1f8" => DATA <= x"05c0";
            when "11" & x"1f9" => DATA <= x"0e07";
            when "11" & x"1fa" => DATA <= x"fbf0";
            when "11" & x"1fb" => DATA <= x"0940";
            when "11" & x"1fc" => DATA <= x"0040";
            when "11" & x"1fd" => DATA <= x"0547";
            when "11" & x"1fe" => DATA <= x"a0ea";
            when "11" & x"1ff" => DATA <= x"0001";
            when "11" & x"200" => DATA <= x"501f";
            when "11" & x"201" => DATA <= x"ffff";
            when "11" & x"202" => DATA <= x"f5fe";
            when "11" & x"203" => DATA <= x"0194";
            when "11" & x"204" => DATA <= x"1a01";
            when "11" & x"205" => DATA <= x"20f9";
            when "11" & x"206" => DATA <= x"b002";
            when "11" & x"207" => DATA <= x"ffc0";
            when "11" & x"208" => DATA <= x"600a";
            when "11" & x"209" => DATA <= x"3feb";
            when "11" & x"20a" => DATA <= x"f008";
            when "11" & x"20b" => DATA <= x"007d";
            when "11" & x"20c" => DATA <= x"c00f";
            when "11" & x"20d" => DATA <= x"f1f8";
            when "11" & x"20e" => DATA <= x"0078";
            when "11" & x"20f" => DATA <= x"fce0";
            when "11" & x"210" => DATA <= x"03f9";
            when "11" & x"211" => DATA <= x"f900";
            when "11" & x"212" => DATA <= x"007f";
            when "11" & x"213" => DATA <= x"b888";
            when "11" & x"214" => DATA <= x"0e06";
            when "11" & x"215" => DATA <= x"0381";
            when "11" & x"216" => DATA <= x"c6e7";
            when "11" & x"217" => DATA <= x"77a7";
            when "11" & x"218" => DATA <= x"e87c";
            when "11" & x"219" => DATA <= x"3c17";
            when "11" & x"21a" => DATA <= x"4f86";
            when "11" & x"21b" => DATA <= x"c3f4";
            when "11" & x"21c" => DATA <= x"8ac4";
            when "11" & x"21d" => DATA <= x"a446";
            when "11" & x"21e" => DATA <= x"2915";
            when "11" & x"21f" => DATA <= x"81f7";
            when "11" & x"220" => DATA <= x"ebf7";
            when "11" & x"221" => DATA <= x"b9dd";
            when "11" & x"222" => DATA <= x"eb5e";
            when "11" & x"223" => DATA <= x"e777";
            when "11" & x"224" => DATA <= x"bbf0";
            when "11" & x"225" => DATA <= x"3cff";
            when "11" & x"226" => DATA <= x"0f00";
            when "11" & x"227" => DATA <= x"120b";
            when "11" & x"228" => DATA <= x"caff";
            when "11" & x"229" => DATA <= x"7838";
            when "11" & x"22a" => DATA <= x"5f0f";
            when "11" & x"22b" => DATA <= x"07f8";
            when "11" & x"22c" => DATA <= x"1cbe";
            when "11" & x"22d" => DATA <= x"ff0b";
            when "11" & x"22e" => DATA <= x"8028";
            when "11" & x"22f" => DATA <= x"05fe";
            when "11" & x"230" => DATA <= x"007e";
            when "11" & x"231" => DATA <= x"bfc0";
            when "11" & x"232" => DATA <= x"0200";
            when "11" & x"233" => DATA <= x"0200";
            when "11" & x"234" => DATA <= x"0e00";
            when "11" & x"235" => DATA <= x"2fbf";
            when "11" & x"236" => DATA <= x"c000";
            when "11" & x"237" => DATA <= x"4000";
            when "11" & x"238" => DATA <= x"15fc";
            when "11" & x"239" => DATA <= x"0ea0";
            when "11" & x"23a" => DATA <= x"f000";
            when "11" & x"23b" => DATA <= x"1280";
            when "11" & x"23c" => DATA <= x"1fe0";
            when "11" & x"23d" => DATA <= x"4a00";
            when "11" & x"23e" => DATA <= x"4050";
            when "11" & x"23f" => DATA <= x"0081";
            when "11" & x"240" => DATA <= x"fe48";
            when "11" & x"241" => DATA <= x"a000";
            when "11" & x"242" => DATA <= x"0d00";
            when "11" & x"243" => DATA <= x"081f";
            when "11" & x"244" => DATA <= x"e02a";
            when "11" & x"245" => DATA <= x"0048";
            when "11" & x"246" => DATA <= x"0810";
            when "11" & x"247" => DATA <= x"0c07";
            when "11" & x"248" => DATA <= x"f9b0";
            when "11" & x"249" => DATA <= x"042f";
            when "11" & x"24a" => DATA <= x"5800";
            when "11" & x"24b" => DATA <= x"5c0f";
            when "11" & x"24c" => DATA <= x"17ed";
            when "11" & x"24d" => DATA <= x"0200";
            when "11" & x"24e" => DATA <= x"c00b";
            when "11" & x"24f" => DATA <= x"f1f9";
            when "11" & x"250" => DATA <= x"fdfe";
            when "11" & x"251" => DATA <= x"0404";
            when "11" & x"252" => DATA <= x"5003";
            when "11" & x"253" => DATA <= x"ec00";
            when "11" & x"254" => DATA <= x"100f";
            when "11" & x"255" => DATA <= x"8207";
            when "11" & x"256" => DATA <= x"4420";
            when "11" & x"257" => DATA <= x"03fc";
            when "11" & x"258" => DATA <= x"0080";
            when "11" & x"259" => DATA <= x"7a00";
            when "11" & x"25a" => DATA <= x"2820";
            when "11" & x"25b" => DATA <= x"00ff";
            when "11" & x"25c" => DATA <= x"402f";
            when "11" & x"25d" => DATA <= x"dff2";
            when "11" & x"25e" => DATA <= x"00ff";
            when "11" & x"25f" => DATA <= x"1800";
            when "11" & x"260" => DATA <= x"1832";
            when "11" & x"261" => DATA <= x"00ff";
            when "11" & x"262" => DATA <= x"a001";
            when "11" & x"263" => DATA <= x"dc80";
            when "11" & x"264" => DATA <= x"3fc4";
            when "11" & x"265" => DATA <= x"4047";
            when "11" & x"266" => DATA <= x"da03";
            when "11" & x"267" => DATA <= x"801b";
            when "11" & x"268" => DATA <= x"f400";
            when "11" & x"269" => DATA <= x"017f";
            when "11" & x"26a" => DATA <= x"f003";
            when "11" & x"26b" => DATA <= x"7e80";
            when "11" & x"26c" => DATA <= x"018f";
            when "11" & x"26d" => DATA <= x"fe00";
            when "11" & x"26e" => DATA <= x"7f90";
            when "11" & x"26f" => DATA <= x"1000";
            when "11" & x"270" => DATA <= x"07f8";
            when "11" & x"271" => DATA <= x"014c";
            when "11" & x"272" => DATA <= x"007f";
            when "11" & x"273" => DATA <= x"8002";
            when "11" & x"274" => DATA <= x"0003";
            when "11" & x"275" => DATA <= x"f800";
            when "11" & x"276" => DATA <= x"1010";
            when "11" & x"277" => DATA <= x"0fb0";
            when "11" & x"278" => DATA <= x"580f";
            when "11" & x"279" => DATA <= x"f56f";
            when "11" & x"27a" => DATA <= x"003f";
            when "11" & x"27b" => DATA <= x"1fe7";
            when "11" & x"27c" => DATA <= x"f67b";
            when "11" & x"27d" => DATA <= x"f380";
            when "11" & x"27e" => DATA <= x"0a65";
            when "11" & x"27f" => DATA <= x"b058";
            when "11" & x"280" => DATA <= x"10fc";
            when "11" & x"281" => DATA <= x"01a0";
            when "11" & x"282" => DATA <= x"007d";
            when "11" & x"283" => DATA <= x"7f88";
            when "11" & x"284" => DATA <= x"0944";
            when "11" & x"285" => DATA <= x"0080";
            when "11" & x"286" => DATA <= x"0130";
            when "11" & x"287" => DATA <= x"6379";
            when "11" & x"288" => DATA <= x"3c00";
            when "11" & x"289" => DATA <= x"2004";
            when "11" & x"28a" => DATA <= x"0000";
            when "11" & x"28b" => DATA <= x"0340";
            when "11" & x"28c" => DATA <= x"0070";
            when "11" & x"28d" => DATA <= x"1800";
            when "11" & x"28e" => DATA <= x"0740";
            when "11" & x"28f" => DATA <= x"0274";
            when "11" & x"290" => DATA <= x"187d";
            when "11" & x"291" => DATA <= x"fe00";
            when "11" & x"292" => DATA <= x"0800";
            when "11" & x"293" => DATA <= x"0102";
            when "11" & x"294" => DATA <= x"5060";
            when "11" & x"295" => DATA <= x"1002";
            when "11" & x"296" => DATA <= x"0464";
            when "11" & x"297" => DATA <= x"8015";
            when "11" & x"298" => DATA <= x"0043";
            when "11" & x"299" => DATA <= x"5021";
            when "11" & x"29a" => DATA <= x"e26c";
            when "11" & x"29b" => DATA <= x"4000";
            when "11" & x"29c" => DATA <= x"0049";
            when "11" & x"29d" => DATA <= x"9a00";
            when "11" & x"29e" => DATA <= x"7fd6";
            when "11" & x"29f" => DATA <= x"f801";
            when "11" & x"2a0" => DATA <= x"ead4";
            when "11" & x"2a1" => DATA <= x"6850";
            when "11" & x"2a2" => DATA <= x"057a";
            when "11" & x"2a3" => DATA <= x"0001";
            when "11" & x"2a4" => DATA <= x"6110";
            when "11" & x"2a5" => DATA <= x"c070";
            when "11" & x"2a6" => DATA <= x"0cf0";
            when "11" & x"2a7" => DATA <= x"0378";
            when "11" & x"2a8" => DATA <= x"0302";
            when "11" & x"2a9" => DATA <= x"800f";
            when "11" & x"2aa" => DATA <= x"80d0";
            when "11" & x"2ab" => DATA <= x"0040";
            when "11" & x"2ac" => DATA <= x"00ff";
            when "11" & x"2ad" => DATA <= x"a001";
            when "11" & x"2ae" => DATA <= x"1500";
            when "11" & x"2af" => DATA <= x"0800";
            when "11" & x"2b0" => DATA <= x"007a";
            when "11" & x"2b1" => DATA <= x"0008";
            when "11" & x"2b2" => DATA <= x"4800";
            when "11" & x"2b3" => DATA <= x"83c0";
            when "11" & x"2b4" => DATA <= x"081e";
            when "11" & x"2b5" => DATA <= x"0054";
            when "11" & x"2b6" => DATA <= x"a004";
            when "11" & x"2b7" => DATA <= x"0480";
            when "11" & x"2b8" => DATA <= x"1068";
            when "11" & x"2b9" => DATA <= x"0081";
            when "11" & x"2ba" => DATA <= x"c004";
            when "11" & x"2bb" => DATA <= x"030d";
            when "11" & x"2bc" => DATA <= x"0000";
            when "11" & x"2bd" => DATA <= x"a800";
            when "11" & x"2be" => DATA <= x"0400";
            when "11" & x"2bf" => DATA <= x"1850";
            when "11" & x"2c0" => DATA <= x"0006";
            when "11" & x"2c1" => DATA <= x"4003";
            when "11" & x"2c2" => DATA <= x"dec0";
            when "11" & x"2c3" => DATA <= x"6af0";
            when "11" & x"2c4" => DATA <= x"0026";
            when "11" & x"2c5" => DATA <= x"8010";
            when "11" & x"2c6" => DATA <= x"0082";
            when "11" & x"2c7" => DATA <= x"07f7";
            when "11" & x"2c8" => DATA <= x"0e27";
            when "11" & x"2c9" => DATA <= x"03c1";
            when "11" & x"2ca" => DATA <= x"a0e3";
            when "11" & x"2cb" => DATA <= x"ff80";
            when "11" & x"2cc" => DATA <= x"03bc";
            when "11" & x"2cd" => DATA <= x"00ff";
            when "11" & x"2ce" => DATA <= x"d000";
            when "11" & x"2cf" => DATA <= x"0801";
            when "11" & x"2d0" => DATA <= x"ffe0";
            when "11" & x"2d1" => DATA <= x"0ffb";
            when "11" & x"2d2" => DATA <= x"0010";
            when "11" & x"2d3" => DATA <= x"bfec";
            when "11" & x"2d4" => DATA <= x"0020";
            when "11" & x"2d5" => DATA <= x"fff0";
            when "11" & x"2d6" => DATA <= x"07ff";
            when "11" & x"2d7" => DATA <= x"0001";
            when "11" & x"2d8" => DATA <= x"3801";
            when "11" & x"2d9" => DATA <= x"fe00";
            when "11" & x"2da" => DATA <= x"4068";
            when "11" & x"2db" => DATA <= x"03fe";
            when "11" & x"2dc" => DATA <= x"4000";
            when "11" & x"2dd" => DATA <= x"5400";
            when "11" & x"2de" => DATA <= x"ffb0";
            when "11" & x"2df" => DATA <= x"0603";
            when "11" & x"2e0" => DATA <= x"fff0";
            when "11" & x"2e1" => DATA <= x"00e2";
            when "11" & x"2e2" => DATA <= x"95d0";
            when "11" & x"2e3" => DATA <= x"e576";
            when "11" & x"2e4" => DATA <= x"2900";
            when "11" & x"2e5" => DATA <= x"aee9";
            when "11" & x"2e6" => DATA <= x"0082";
            when "11" & x"2e7" => DATA <= x"4002";
            when "11" & x"2e8" => DATA <= x"d000";
            when "11" & x"2e9" => DATA <= x"5c28";
            when "11" & x"2ea" => DATA <= x"806b";
            when "11" & x"2eb" => DATA <= x"2000";
            when "11" & x"2ec" => DATA <= x"0d57";
            when "11" & x"2ed" => DATA <= x"ab55";
            when "11" & x"2ee" => DATA <= x"51d5";
            when "11" & x"2ef" => DATA <= x"2a85";
            when "11" & x"2f0" => DATA <= x"7aad";
            when "11" & x"2f1" => DATA <= x"9f50";
            when "11" & x"2f2" => DATA <= x"0835";
            when "11" & x"2f3" => DATA <= x"8a8d";
            when "11" & x"2f4" => DATA <= x"e6a7";
            when "11" & x"2f5" => DATA <= x"4597";
            when "11" & x"2f6" => DATA <= x"edfc";
            when "11" & x"2f7" => DATA <= x"8f40";
            when "11" & x"2f8" => DATA <= x"0c56";
            when "11" & x"2f9" => DATA <= x"0821";
            when "11" & x"2fa" => DATA <= x"f8f8";
            when "11" & x"2fb" => DATA <= x"0036";
            when "11" & x"2fc" => DATA <= x"1f8f";
            when "11" & x"2fd" => DATA <= x"f008";
            when "11" & x"2fe" => DATA <= x"02bf";
            when "11" & x"2ff" => DATA <= x"c000";
            when "11" & x"300" => DATA <= x"4408";
            when "11" & x"301" => DATA <= x"3e80";
            when "11" & x"302" => DATA <= x"2bfd";
            when "11" & x"303" => DATA <= x"c15f";
            when "11" & x"304" => DATA <= x"eefa";
            when "11" & x"305" => DATA <= x"005f";
            when "11" & x"306" => DATA <= x"effb";
            when "11" & x"307" => DATA <= x"e9f9";
            when "11" & x"308" => DATA <= x"dfe4";
            when "11" & x"309" => DATA <= x"1f01";
            when "11" & x"30a" => DATA <= x"f000";
            when "11" & x"30b" => DATA <= x"03c3";
            when "11" & x"30c" => DATA <= x"ffc7";
            when "11" & x"30d" => DATA <= x"e2fb";
            when "11" & x"30e" => DATA <= x"3fb0";
            when "11" & x"30f" => DATA <= x"0afc";
            when "11" & x"310" => DATA <= x"b00a";
            when "11" & x"311" => DATA <= x"ff73";
            when "11" & x"312" => DATA <= x"002b";
            when "11" & x"313" => DATA <= x"8080";
            when "11" & x"314" => DATA <= x"e667";
            when "11" & x"315" => DATA <= x"b1d3";
            when "11" & x"316" => DATA <= x"f43e";
            when "11" & x"317" => DATA <= x"9f0f";
            when "11" & x"318" => DATA <= x"a7c3";
            when "11" & x"319" => DATA <= x"e1b6";
            when "11" & x"31a" => DATA <= x"2314";
            when "11" & x"31b" => DATA <= x"0a45";
            when "11" & x"31c" => DATA <= x"20d2";
            when "11" & x"31d" => DATA <= x"0110";
            when "11" & x"31e" => DATA <= x"ff57";
            when "11" & x"31f" => DATA <= x"f4ff";
            when "11" & x"320" => DATA <= x"dfe3";
            when "11" & x"321" => DATA <= x"ca37";
            when "11" & x"322" => DATA <= x"0c1f";
            when "11" & x"323" => DATA <= x"1c60";
            when "11" & x"324" => DATA <= x"7428";
            when "11" & x"325" => DATA <= x"b380";
            when "11" & x"326" => DATA <= x"090b";
            when "11" & x"327" => DATA <= x"7401";
            when "11" & x"328" => DATA <= x"041e";
            when "11" & x"329" => DATA <= x"0008";
            when "11" & x"32a" => DATA <= x"0004";
            when "11" & x"32b" => DATA <= x"8f70";
            when "11" & x"32c" => DATA <= x"2001";
            when "11" & x"32d" => DATA <= x"fef8";
            when "11" & x"32e" => DATA <= x"7e34";
            when "11" & x"32f" => DATA <= x"1060";
            when "11" & x"330" => DATA <= x"6430";
            when "11" & x"331" => DATA <= x"027f";
            when "11" & x"332" => DATA <= x"c3c0";
            when "11" & x"333" => DATA <= x"0010";
            when "11" & x"334" => DATA <= x"002e";
            when "11" & x"335" => DATA <= x"02e1";
            when "11" & x"336" => DATA <= x"f000";
            when "11" & x"337" => DATA <= x"7838";
            when "11" & x"338" => DATA <= x"1000";
            when "11" & x"339" => DATA <= x"0104";
            when "11" & x"33a" => DATA <= x"1e00";
            when "11" & x"33b" => DATA <= x"f010";
            when "11" & x"33c" => DATA <= x"8040";
            when "11" & x"33d" => DATA <= x"6b80";
            when "11" & x"33e" => DATA <= x"03fc";
            when "11" & x"33f" => DATA <= x"00ff";
            when "11" & x"340" => DATA <= x"2204";
            when "11" & x"341" => DATA <= x"4021";
            when "11" & x"342" => DATA <= x"1101";
            when "11" & x"343" => DATA <= x"fc00";
            when "11" & x"344" => DATA <= x"7e04";
            when "11" & x"345" => DATA <= x"0880";
            when "11" & x"346" => DATA <= x"4c30";
            when "11" & x"347" => DATA <= x"80d0";
            when "11" & x"348" => DATA <= x"00f4";
            when "11" & x"349" => DATA <= x"e000";
            when "11" & x"34a" => DATA <= x"1002";
            when "11" & x"34b" => DATA <= x"805f";
            when "11" & x"34c" => DATA <= x"bc00";
            when "11" & x"34d" => DATA <= x"0300";
            when "11" & x"34e" => DATA <= x"9040";
            when "11" & x"34f" => DATA <= x"0ffa";
            when "11" & x"350" => DATA <= x"0008";
            when "11" & x"351" => DATA <= x"0481";
            when "11" & x"352" => DATA <= x"8b87";
            when "11" & x"353" => DATA <= x"600e";
            when "11" & x"354" => DATA <= x"8000";
            when "11" & x"355" => DATA <= x"4120";
            when "11" & x"356" => DATA <= x"231c";
            when "11" & x"357" => DATA <= x"4c08";
            when "11" & x"358" => DATA <= x"e000";
            when "11" & x"359" => DATA <= x"4000";
            when "11" & x"35a" => DATA <= x"88f0";
            when "11" & x"35b" => DATA <= x"0810";
            when "11" & x"35c" => DATA <= x"0015";
            when "11" & x"35d" => DATA <= x"0140";
            when "11" & x"35e" => DATA <= x"0fa2";
            when "11" & x"35f" => DATA <= x"03e0";
            when "11" & x"360" => DATA <= x"00f0";
            when "11" & x"361" => DATA <= x"e005";
            when "11" & x"362" => DATA <= x"5808";
            when "11" & x"363" => DATA <= x"0200";
            when "11" & x"364" => DATA <= x"7fa3";
            when "11" & x"365" => DATA <= x"2801";
            when "11" & x"366" => DATA <= x"fe00";
            when "11" & x"367" => DATA <= x"100d";
            when "11" & x"368" => DATA <= x"100e";
            when "11" & x"369" => DATA <= x"6101";
            when "11" & x"36a" => DATA <= x"a1f2";
            when "11" & x"36b" => DATA <= x"0062";
            when "11" & x"36c" => DATA <= x"3440";
            when "11" & x"36d" => DATA <= x"2627";
            when "11" & x"36e" => DATA <= x"c001";
            when "11" & x"36f" => DATA <= x"fe00";
            when "11" & x"370" => DATA <= x"00af";
            when "11" & x"371" => DATA <= x"6800";
            when "11" & x"372" => DATA <= x"0208";
            when "11" & x"373" => DATA <= x"7f80";
            when "11" & x"374" => DATA <= x"0408";
            when "11" & x"375" => DATA <= x"0000";
            when "11" & x"376" => DATA <= x"4280";
            when "11" & x"377" => DATA <= x"1fe0";
            when "11" & x"378" => DATA <= x"0008";
            when "11" & x"379" => DATA <= x"9240";
            when "11" & x"37a" => DATA <= x"1fe0";
            when "11" & x"37b" => DATA <= x"0008";
            when "11" & x"37c" => DATA <= x"4421";
            when "11" & x"37d" => DATA <= x"c00f";
            when "11" & x"37e" => DATA <= x"f782";
            when "11" & x"37f" => DATA <= x"c288";
            when "11" & x"380" => DATA <= x"3800";
            when "11" & x"381" => DATA <= x"2201";
            when "11" & x"382" => DATA <= x"7b82";
            when "11" & x"383" => DATA <= x"6801";
            when "11" & x"384" => DATA <= x"00bc";
            when "11" & x"385" => DATA <= x"5fa0";
            when "11" & x"386" => DATA <= x"1fef";
            when "11" & x"387" => DATA <= x"ba18";
            when "11" & x"388" => DATA <= x"9030";
            when "11" & x"389" => DATA <= x"3bbe";
            when "11" & x"38a" => DATA <= x"4018";
            when "11" & x"38b" => DATA <= x"0206";
            when "11" & x"38c" => DATA <= x"e3f6";
            when "11" & x"38d" => DATA <= x"8000";
            when "11" & x"38e" => DATA <= x"2c00";
            when "11" & x"38f" => DATA <= x"287c";
            when "11" & x"390" => DATA <= x"aef7";
            when "11" & x"391" => DATA <= x"138d";
            when "11" & x"392" => DATA <= x"6401";
            when "11" & x"393" => DATA <= x"9cff";
            when "11" & x"394" => DATA <= x"0703";
            when "11" & x"395" => DATA <= x"2b7d";
            when "11" & x"396" => DATA <= x"80d0";
            when "11" & x"397" => DATA <= x"aff7";
            when "11" & x"398" => DATA <= x"b111";
            when "11" & x"399" => DATA <= x"e8fc";
            when "11" & x"39a" => DATA <= x"024f";
            when "11" & x"39b" => DATA <= x"f8d1";
            when "11" & x"39c" => DATA <= x"1ccf";
            when "11" & x"39d" => DATA <= x"0057";
            when "11" & x"39e" => DATA <= x"fa7c";
            when "11" & x"39f" => DATA <= x"1a00";
            when "11" & x"3a0" => DATA <= x"783f";
            when "11" & x"3a1" => DATA <= x"c015";
            when "11" & x"3a2" => DATA <= x"fe1f";
            when "11" & x"3a3" => DATA <= x"0008";
            when "11" & x"3a4" => DATA <= x"abfc";
            when "11" & x"3a5" => DATA <= x"015f";
            when "11" & x"3a6" => DATA <= x"ec04";
            when "11" & x"3a7" => DATA <= x"0304";
            when "11" & x"3a8" => DATA <= x"868f";
            when "11" & x"3a9" => DATA <= x"003f";
            when "11" & x"3aa" => DATA <= x"e47c";
            when "11" & x"3ab" => DATA <= x"1000";
            when "11" & x"3ac" => DATA <= x"083f";
            when "11" & x"3ad" => DATA <= x"f400";
            when "11" & x"3ae" => DATA <= x"0400";
            when "11" & x"3af" => DATA <= x"7fc8";
            when "11" & x"3b0" => DATA <= x"0281";
            when "11" & x"3b1" => DATA <= x"5201";
            when "11" & x"3b2" => DATA <= x"7f80";
            when "11" & x"3b3" => DATA <= x"f806";
            when "11" & x"3b4" => DATA <= x"a284";
            when "11" & x"3b5" => DATA <= x"0ff1";
            when "11" & x"3b6" => DATA <= x"8710";
            when "11" & x"3b7" => DATA <= x"2108";
            when "11" & x"3b8" => DATA <= x"4007";
            when "11" & x"3b9" => DATA <= x"fc80";
            when "11" & x"3ba" => DATA <= x"280a";
            when "11" & x"3bb" => DATA <= x"2027";
            when "11" & x"3bc" => DATA <= x"ff03";
            when "11" & x"3bd" => DATA <= x"0081";
            when "11" & x"3be" => DATA <= x"4050";
            when "11" & x"3bf" => DATA <= x"03fe";
            when "11" & x"3c0" => DATA <= x"400c";
            when "11" & x"3c1" => DATA <= x"06a3";
            when "11" & x"3c2" => DATA <= x"41fc";
            when "11" & x"3c3" => DATA <= x"614e";
            when "11" & x"3c4" => DATA <= x"0740";
            when "11" & x"3c5" => DATA <= x"2d00";
            when "11" & x"3c6" => DATA <= x"0428";
            when "11" & x"3c7" => DATA <= x"0009";
            when "11" & x"3c8" => DATA <= x"2000";
            when "11" & x"3c9" => DATA <= x"c200";
            when "11" & x"3ca" => DATA <= x"0140";
            when "11" & x"3cb" => DATA <= x"c00f";
            when "11" & x"3cc" => DATA <= x"50e1";
            when "11" & x"3cd" => DATA <= x"783c";
            when "11" & x"3ce" => DATA <= x"3c0e";
            when "11" & x"3cf" => DATA <= x"07e8";
            when "11" & x"3d0" => DATA <= x"0022";
            when "11" & x"3d1" => DATA <= x"1000";
            when "11" & x"3d2" => DATA <= x"0400";
            when "11" & x"3d3" => DATA <= x"5200";
            when "11" & x"3d4" => DATA <= x"11b0";
            when "11" & x"3d5" => DATA <= x"0400";
            when "11" & x"3d6" => DATA <= x"2800";
            when "11" & x"3d7" => DATA <= x"80a0";
            when "11" & x"3d8" => DATA <= x"0082";
            when "11" & x"3d9" => DATA <= x"0005";
            when "11" & x"3da" => DATA <= x"6000";
            when "11" & x"3db" => DATA <= x"1061";
            when "11" & x"3dc" => DATA <= x"4280";
            when "11" & x"3dd" => DATA <= x"021c";
            when "11" & x"3de" => DATA <= x"0002";
            when "11" & x"3df" => DATA <= x"3070";
            when "11" & x"3e0" => DATA <= x"0200";
            when "11" & x"3e1" => DATA <= x"3024";
            when "11" & x"3e2" => DATA <= x"e000";
            when "11" & x"3e3" => DATA <= x"1480";
            when "11" & x"3e4" => DATA <= x"182c";
            when "11" & x"3e5" => DATA <= x"0004";
            when "11" & x"3e6" => DATA <= x"fc02";
            when "11" & x"3e7" => DATA <= x"3480";
            when "11" & x"3e8" => DATA <= x"042e";
            when "11" & x"3e9" => DATA <= x"0046";
            when "11" & x"3ea" => DATA <= x"8012";
            when "11" & x"3eb" => DATA <= x"c001";
            when "11" & x"3ec" => DATA <= x"1500";
            when "11" & x"3ed" => DATA <= x"1009";
            when "11" & x"3ee" => DATA <= x"8004";
            when "11" & x"3ef" => DATA <= x"b000";
            when "11" & x"3f0" => DATA <= x"2400";
            when "11" & x"3f1" => DATA <= x"1d2e";
            when "11" & x"3f2" => DATA <= x"a8e9";
            when "11" & x"3f3" => DATA <= x"743a";
            when "11" & x"3f4" => DATA <= x"1d8e";
            when "11" & x"3f5" => DATA <= x"801e";
            when "11" & x"3f6" => DATA <= x"abfa";
            when "11" & x"3f7" => DATA <= x"ad59";
            when "11" & x"3f8" => DATA <= x"ab9a";
            when "11" & x"3f9" => DATA <= x"9552";
            when "11" & x"3fa" => DATA <= x"b516";
            when "11" & x"3fb" => DATA <= x"8175";
            when "11" & x"3fc" => DATA <= x"3ad5";
            when "11" & x"3fd" => DATA <= x"4ea3";
            when "11" & x"3fe" => DATA <= x"f9bd";
            when "11" & x"3ff" => DATA <= x"fe5f";
            when "11" & x"400" => DATA <= x"3fbd";
            when "11" & x"401" => DATA <= x"e9fc";
            when "11" & x"402" => DATA <= x"2000";
            when "11" & x"403" => DATA <= x"7c80";
            when "11" & x"404" => DATA <= x"0100";
            when "11" & x"405" => DATA <= x"27e3";
            when "11" & x"406" => DATA <= x"e280";
            when "11" & x"407" => DATA <= x"007c";
            when "11" & x"408" => DATA <= x"00ff";
            when "11" & x"409" => DATA <= x"07a0";
            when "11" & x"40a" => DATA <= x"0015";
            when "11" & x"40b" => DATA <= x"00c0";
            when "11" & x"40c" => DATA <= x"703f";
            when "11" & x"40d" => DATA <= x"c1ff";
            when "11" & x"40e" => DATA <= x"fe00";
            when "11" & x"40f" => DATA <= x"fff7";
            when "11" & x"410" => DATA <= x"b500";
            when "11" & x"411" => DATA <= x"9c74";
            when "11" & x"412" => DATA <= x"07c0";
            when "11" & x"413" => DATA <= x"0015";
            when "11" & x"414" => DATA <= x"fe07";
            when "11" & x"415" => DATA <= x"0030";
            when "11" & x"416" => DATA <= x"1f95";
            when "11" & x"417" => DATA <= x"fe3f";
            when "11" & x"418" => DATA <= x"0020";
            when "11" & x"419" => DATA <= x"1795";
            when "11" & x"41a" => DATA <= x"7e3f";
            when "11" & x"41b" => DATA <= x"5fd0";
            when "11" & x"41c" => DATA <= x"03ff";
            when "11" & x"41d" => DATA <= x"c00f";
            when "11" & x"41e" => DATA <= x"fa00";
            when "11" & x"41f" => DATA <= x"e7ee";
            when "11" & x"420" => DATA <= x"0005";
            when "11" & x"421" => DATA <= x"7130";
            when "11" & x"422" => DATA <= x"13e1";
            when "11" & x"423" => DATA <= x"f0f7";
            when "11" & x"424" => DATA <= x"0fa7";
            when "11" & x"425" => DATA <= x"c3e4";
            when "11" & x"426" => DATA <= x"5a44";
            when "11" & x"427" => DATA <= x"2011";
            when "11" & x"428" => DATA <= x"6934";
            when "11" & x"429" => DATA <= x"0b5f";
            when "11" & x"42a" => DATA <= x"f2fe";
            when "11" & x"42b" => DATA <= x"7e3f";
            when "11" & x"42c" => DATA <= x"f009";
            when "11" & x"42d" => DATA <= x"cd26";
            when "11" & x"42e" => DATA <= x"c329";
            when "11" & x"42f" => DATA <= x"9ec4";
            when "11" & x"430" => DATA <= x"1480";
            when "11" & x"431" => DATA <= x"912c";
            when "11" & x"432" => DATA <= x"1918";
            when "11" & x"433" => DATA <= x"0000";
            when "11" & x"434" => DATA <= x"1500";
            when "11" & x"435" => DATA <= x"3dc8";
            when "11" & x"436" => DATA <= x"4020";
            when "11" & x"437" => DATA <= x"2023";
            when "11" & x"438" => DATA <= x"801f";
            when "11" & x"439" => DATA <= x"ede1";
            when "11" & x"43a" => DATA <= x"0000";
            when "11" & x"43b" => DATA <= x"1140";
            when "11" & x"43c" => DATA <= x"0087";
            when "11" & x"43d" => DATA <= x"f800";
            when "11" & x"43e" => DATA <= x"0209";
            when "11" & x"43f" => DATA <= x"1087";
            when "11" & x"440" => DATA <= x"0e08";
            when "11" & x"441" => DATA <= x"a25a";
            when "11" & x"442" => DATA <= x"91c8";
            when "11" & x"443" => DATA <= x"05e0";
            when "11" & x"444" => DATA <= x"009a";
            when "11" & x"445" => DATA <= x"71c6";
            when "11" & x"446" => DATA <= x"011f";
            when "11" & x"447" => DATA <= x"3803";
            when "11" & x"448" => DATA <= x"080a";
            when "11" & x"449" => DATA <= x"00af";
            when "11" & x"44a" => DATA <= x"f3f8";
            when "11" & x"44b" => DATA <= x"6000";
            when "11" & x"44c" => DATA <= x"f7a0";
            when "11" & x"44d" => DATA <= x"0aff";
            when "11" & x"44e" => DATA <= x"e007";
            when "11" & x"44f" => DATA <= x"bd00";
            when "11" & x"450" => DATA <= x"57ff";
            when "11" & x"451" => DATA <= x"003f";
            when "11" & x"452" => DATA <= x"e800";
            when "11" & x"453" => DATA <= x"3eff";
            when "11" & x"454" => DATA <= x"6614";
            when "11" & x"455" => DATA <= x"1000";
            when "11" & x"456" => DATA <= x"e36b";
            when "11" & x"457" => DATA <= x"8100";
            when "11" & x"458" => DATA <= x"0000";
            when "11" & x"459" => DATA <= x"8ec3";
            when "11" & x"45a" => DATA <= x"e782";
            when "11" & x"45b" => DATA <= x"c02c";
            when "11" & x"45c" => DATA <= x"6214";
            when "11" & x"45d" => DATA <= x"6000";
            when "11" & x"45e" => DATA <= x"0049";
            when "11" & x"45f" => DATA <= x"2090";
            when "11" & x"460" => DATA <= x"1cc4";
            when "11" & x"461" => DATA <= x"667f";
            when "11" & x"462" => DATA <= x"bf81";
            when "11" & x"463" => DATA <= x"04d0";
            when "11" & x"464" => DATA <= x"0831";
            when "11" & x"465" => DATA <= x"1880";
            when "11" & x"466" => DATA <= x"0302";
            when "11" & x"467" => DATA <= x"1015";
            when "11" & x"468" => DATA <= x"8087";
            when "11" & x"469" => DATA <= x"4b8b";
            when "11" & x"46a" => DATA <= x"df80";
            when "11" & x"46b" => DATA <= x"00f0";
            when "11" & x"46c" => DATA <= x"01e0";
            when "11" & x"46d" => DATA <= x"000f";
            when "11" & x"46e" => DATA <= x"801f";
            when "11" & x"46f" => DATA <= x"e000";
            when "11" & x"470" => DATA <= x"6230";
            when "11" & x"471" => DATA <= x"1f5f";
            when "11" & x"472" => DATA <= x"85c1";
            when "11" & x"473" => DATA <= x"fd00";
            when "11" & x"474" => DATA <= x"5603";
            when "11" & x"475" => DATA <= x"1c02";
            when "11" & x"476" => DATA <= x"8007";
            when "11" & x"477" => DATA <= x"7002";
            when "11" & x"478" => DATA <= x"812c";
            when "11" & x"479" => DATA <= x"0103";
            when "11" & x"47a" => DATA <= x"1010";
            when "11" & x"47b" => DATA <= x"000a";
            when "11" & x"47c" => DATA <= x"405b";
            when "11" & x"47d" => DATA <= x"a103";
            when "11" & x"47e" => DATA <= x"0010";
            when "11" & x"47f" => DATA <= x"9000";
            when "11" & x"480" => DATA <= x"1800";
            when "11" & x"481" => DATA <= x"7f85";
            when "11" & x"482" => DATA <= x"8a1c";
            when "11" & x"483" => DATA <= x"0040";
            when "11" & x"484" => DATA <= x"001f";
            when "11" & x"485" => DATA <= x"d834";
            when "11" & x"486" => DATA <= x"0009";
            when "11" & x"487" => DATA <= x"e003";
            when "11" & x"488" => DATA <= x"e001";
            when "11" & x"489" => DATA <= x"0481";
            when "11" & x"48a" => DATA <= x"4150";
            when "11" & x"48b" => DATA <= x"01f9";
            when "11" & x"48c" => DATA <= x"8000";
            when "11" & x"48d" => DATA <= x"6010";
            when "11" & x"48e" => DATA <= x"041c";
            when "11" & x"48f" => DATA <= x"0080";
            when "11" & x"490" => DATA <= x"a40a";
            when "11" & x"491" => DATA <= x"c0a0";
            when "11" & x"492" => DATA <= x"8025";
            when "11" & x"493" => DATA <= x"00f8";
            when "11" & x"494" => DATA <= x"0680";
            when "11" & x"495" => DATA <= x"0a29";
            when "11" & x"496" => DATA <= x"0011";
            when "11" & x"497" => DATA <= x"4008";
            when "11" & x"498" => DATA <= x"0001";
            when "11" & x"499" => DATA <= x"0000";
            when "11" & x"49a" => DATA <= x"2504";
            when "11" & x"49b" => DATA <= x"5091";
            when "11" & x"49c" => DATA <= x"8800";
            when "11" & x"49d" => DATA <= x"0d4c";
            when "11" & x"49e" => DATA <= x"0000";
            when "11" & x"49f" => DATA <= x"5400";
            when "11" & x"4a0" => DATA <= x"1800";
            when "11" & x"4a1" => DATA <= x"1028";
            when "11" & x"4a2" => DATA <= x"0011";
            when "11" & x"4a3" => DATA <= x"4001";
            when "11" & x"4a4" => DATA <= x"8001";
            when "11" & x"4a5" => DATA <= x"4802";
            when "11" & x"4a6" => DATA <= x"0030";
            when "11" & x"4a7" => DATA <= x"0000";
            when "11" & x"4a8" => DATA <= x"4080";
            when "11" & x"4a9" => DATA <= x"0014";
            when "11" & x"4aa" => DATA <= x"10d0";
            when "11" & x"4ab" => DATA <= x"6701";
            when "11" & x"4ac" => DATA <= x"2800";
            when "11" & x"4ad" => DATA <= x"0408";
            when "11" & x"4ae" => DATA <= x"5829";
            when "11" & x"4af" => DATA <= x"122a";
            when "11" & x"4b0" => DATA <= x"8640";
            when "11" & x"4b1" => DATA <= x"02bc";
            when "11" & x"4b2" => DATA <= x"3bfd";
            when "11" & x"4b3" => DATA <= x"c0c0";
            when "11" & x"4b4" => DATA <= x"0170";
            when "11" & x"4b5" => DATA <= x"f83c";
            when "11" & x"4b6" => DATA <= x"3e0f";
            when "11" & x"4b7" => DATA <= x"7f80";
            when "11" & x"4b8" => DATA <= x"121a";
            when "11" & x"4b9" => DATA <= x"003f";
            when "11" & x"4ba" => DATA <= x"1c02";
            when "11" & x"4bb" => DATA <= x"bc00";
            when "11" & x"4bc" => DATA <= x"0200";
            when "11" & x"4bd" => DATA <= x"00e8";
            when "11" & x"4be" => DATA <= x"00c0";
            when "11" & x"4bf" => DATA <= x"0020";
            when "11" & x"4c0" => DATA <= x"f00b";
            when "11" & x"4c1" => DATA <= x"0003";
            when "11" & x"4c2" => DATA <= x"0000";
            when "11" & x"4c3" => DATA <= x"8f04";
            when "11" & x"4c4" => DATA <= x"8143";
            when "11" & x"4c5" => DATA <= x"4028";
            when "11" & x"4c6" => DATA <= x"0c00";
            when "11" & x"4c7" => DATA <= x"027f";
            when "11" & x"4c8" => DATA <= x"1c69";
            when "11" & x"4c9" => DATA <= x"c000";
            when "11" & x"4ca" => DATA <= x"e0a0";
            when "11" & x"4cb" => DATA <= x"07fd";
            when "11" & x"4cc" => DATA <= x"0010";
            when "11" & x"4cd" => DATA <= x"1c0b";
            when "11" & x"4ce" => DATA <= x"7700";
            when "11" & x"4cf" => DATA <= x"01fe";
            when "11" & x"4d0" => DATA <= x"086c";
            when "11" & x"4d1" => DATA <= x"aa5f";
            when "11" & x"4d2" => DATA <= x"c061";
            when "11" & x"4d3" => DATA <= x"f861";
            when "11" & x"4d4" => DATA <= x"fe1c";
            when "11" & x"4d5" => DATA <= x"e1f3";
            when "11" & x"4d6" => DATA <= x"e074";
            when "11" & x"4d7" => DATA <= x"3c1f";
            when "11" & x"4d8" => DATA <= x"a000";
            when "11" & x"4d9" => DATA <= x"1000";
            when "11" & x"4da" => DATA <= x"91a0";
            when "11" & x"4db" => DATA <= x"0420";
            when "11" & x"4dc" => DATA <= x"0203";
            when "11" & x"4dd" => DATA <= x"c02c";
            when "11" & x"4de" => DATA <= x"0012";
            when "11" & x"4df" => DATA <= x"0023";
            when "11" & x"4e0" => DATA <= x"0424";
            when "11" & x"4e1" => DATA <= x"0006";
            when "11" & x"4e2" => DATA <= x"0840";
            when "11" & x"4e3" => DATA <= x"d000";
            when "11" & x"4e4" => DATA <= x"9070";
            when "11" & x"4e5" => DATA <= x"0003";
            when "11" & x"4e6" => DATA <= x"040a";
            when "11" & x"4e7" => DATA <= x"0000";
            when "11" & x"4e8" => DATA <= x"880c";
            when "11" & x"4e9" => DATA <= x"10c0";
            when "11" & x"4ea" => DATA <= x"a004";
            when "11" & x"4eb" => DATA <= x"8001";
            when "11" & x"4ec" => DATA <= x"8140";
            when "11" & x"4ed" => DATA <= x"0294";
            when "11" & x"4ee" => DATA <= x"0000";
            when "11" & x"4ef" => DATA <= x"4003";
            when "11" & x"4f0" => DATA <= x"0e3b";
            when "11" & x"4f1" => DATA <= x"0001";
            when "11" & x"4f2" => DATA <= x"1d00";
            when "11" & x"4f3" => DATA <= x"0380";
            when "11" & x"4f4" => DATA <= x"1412";
            when "11" & x"4f5" => DATA <= x"0004";
            when "11" & x"4f6" => DATA <= x"9006";
            when "11" & x"4f7" => DATA <= x"0391";
            when "11" & x"4f8" => DATA <= x"48e2";
            when "11" & x"4f9" => DATA <= x"602e";
            when "11" & x"4fa" => DATA <= x"aaed";
            when "11" & x"4fb" => DATA <= x"7b5d";
            when "11" & x"4fc" => DATA <= x"d4dd";
            when "11" & x"4fd" => DATA <= x"2aa5";
            when "11" & x"4fe" => DATA <= x"77ed";
            when "11" & x"4ff" => DATA <= x"2ab5";
            when "11" & x"500" => DATA <= x"52ad";
            when "11" & x"501" => DATA <= x"54ad";
            when "11" & x"502" => DATA <= x"6aaf";
            when "11" & x"503" => DATA <= x"deaa";
            when "11" & x"504" => DATA <= x"957c";
            when "11" & x"505" => DATA <= x"d5aa";
            when "11" & x"506" => DATA <= x"5755";
            when "11" & x"507" => DATA <= x"5482";
            when "11" & x"508" => DATA <= x"40d5";
            when "11" & x"509" => DATA <= x"5229";
            when "11" & x"50a" => DATA <= x"1677";
            when "11" & x"50b" => DATA <= x"f7f0";
            when "11" & x"50c" => DATA <= x"0205";
            when "11" & x"50d" => DATA <= x"8b40";
            when "11" & x"50e" => DATA <= x"002e";
            when "11" & x"50f" => DATA <= x"0040";
            when "11" & x"510" => DATA <= x"3fdf";
            when "11" & x"511" => DATA <= x"804a";
            when "11" & x"512" => DATA <= x"0002";
            when "11" & x"513" => DATA <= x"0001";
            when "11" & x"514" => DATA <= x"e8f4";
            when "11" & x"515" => DATA <= x"1d40";
            when "11" & x"516" => DATA <= x"0010";
            when "11" & x"517" => DATA <= x"0e00";
            when "11" & x"518" => DATA <= x"07ff";
            when "11" & x"519" => DATA <= x"b82f";
            when "11" & x"51a" => DATA <= x"ffc0";
            when "11" & x"51b" => DATA <= x"403e";
            when "11" & x"51c" => DATA <= x"0000";
            when "11" & x"51d" => DATA <= x"dff0";
            when "11" & x"51e" => DATA <= x"3800";
            when "11" & x"51f" => DATA <= x"09d7";
            when "11" & x"520" => DATA <= x"e3f0";
            when "11" & x"521" => DATA <= x"0800";
            when "11" & x"522" => DATA <= x"603e";
            when "11" & x"523" => DATA <= x"003f";
            when "11" & x"524" => DATA <= x"cff4";
            when "11" & x"525" => DATA <= x"00fc";
            when "11" & x"526" => DATA <= x"e003";
            when "11" & x"527" => DATA <= x"fbe0";
            when "11" & x"528" => DATA <= x"00fc";
            when "11" & x"529" => DATA <= x"7fd0";
            when "11" & x"52a" => DATA <= x"0560";
            when "11" & x"52b" => DATA <= x"381c";
            when "11" & x"52c" => DATA <= x"6e76";
            when "11" & x"52d" => DATA <= x"7b98";
            when "11" & x"52e" => DATA <= x"001f";
            when "11" & x"52f" => DATA <= x"0f05";
            when "11" & x"530" => DATA <= x"d3e1";
            when "11" & x"531" => DATA <= x"b0fa";
            when "11" & x"532" => DATA <= x"7c3c";
            when "11" & x"533" => DATA <= x"4423";
            when "11" & x"534" => DATA <= x"7229";
            when "11" & x"535" => DATA <= x"0088";
            when "11" & x"536" => DATA <= x"45f7";
            when "11" & x"537" => DATA <= x"f3e9";
            when "11" & x"538" => DATA <= x"ce8c";
            when "11" & x"539" => DATA <= x"d67c";
            when "11" & x"53a" => DATA <= x"a6d3";
            when "11" & x"53b" => DATA <= x"001c";
            when "11" & x"53c" => DATA <= x"000e";
            when "11" & x"53d" => DATA <= x"b09d";
            when "11" & x"53e" => DATA <= x"0080";
            when "11" & x"53f" => DATA <= x"0640";
            when "11" & x"540" => DATA <= x"1000";
            when "11" & x"541" => DATA <= x"3e80";
            when "11" & x"542" => DATA <= x"1000";
            when "11" & x"543" => DATA <= x"02b5";
            when "11" & x"544" => DATA <= x"0020";
            when "11" & x"545" => DATA <= x"2800";
            when "11" & x"546" => DATA <= x"8000";
            when "11" & x"547" => DATA <= x"193f";
            when "11" & x"548" => DATA <= x"8026";
            when "11" & x"549" => DATA <= x"1070";
            when "11" & x"54a" => DATA <= x"0041";
            when "11" & x"54b" => DATA <= x"4000";
            when "11" & x"54c" => DATA <= x"f7e1";
            when "11" & x"54d" => DATA <= x"8418";
            when "11" & x"54e" => DATA <= x"0018";
            when "11" & x"54f" => DATA <= x"5003";
            when "11" & x"550" => DATA <= x"f07e";
            when "11" & x"551" => DATA <= x"3001";
            when "11" & x"552" => DATA <= x"8002";
            when "11" & x"553" => DATA <= x"1400";
            when "11" & x"554" => DATA <= x"2b00";
            when "11" & x"555" => DATA <= x"0f3c";
            when "11" & x"556" => DATA <= x"0000";
            when "11" & x"557" => DATA <= x"0840";
            when "11" & x"558" => DATA <= x"7800";
            when "11" & x"559" => DATA <= x"0100";
            when "11" & x"55a" => DATA <= x"0840";
            when "11" & x"55b" => DATA <= x"0084";
            when "11" & x"55c" => DATA <= x"0040";
            when "11" & x"55d" => DATA <= x"9822";
            when "11" & x"55e" => DATA <= x"a25b";
            when "11" & x"55f" => DATA <= x"440a";
            when "11" & x"560" => DATA <= x"c064";
            when "11" & x"561" => DATA <= x"3380";
            when "11" & x"562" => DATA <= x"6470";
            when "11" & x"563" => DATA <= x"0018";
            when "11" & x"564" => DATA <= x"661f";
            when "11" & x"565" => DATA <= x"aff0";
            when "11" & x"566" => DATA <= x"00a2";
            when "11" & x"567" => DATA <= x"402b";
            when "11" & x"568" => DATA <= x"fd00";
            when "11" & x"569" => DATA <= x"de7c";
            when "11" & x"56a" => DATA <= x"7003";
            when "11" & x"56b" => DATA <= x"fc02";
            when "11" & x"56c" => DATA <= x"c13f";
            when "11" & x"56d" => DATA <= x"f000";
            when "11" & x"56e" => DATA <= x"2d32";
            when "11" & x"56f" => DATA <= x"010f";
            when "11" & x"570" => DATA <= x"8528";
            when "11" & x"571" => DATA <= x"003c";
            when "11" & x"572" => DATA <= x"0000";
            when "11" & x"573" => DATA <= x"851f";
            when "11" & x"574" => DATA <= x"c90a";
            when "11" & x"575" => DATA <= x"007e";
            when "11" & x"576" => DATA <= x"802a";
            when "11" & x"577" => DATA <= x"01a2";
            when "11" & x"578" => DATA <= x"ff40";
            when "11" & x"579" => DATA <= x"0001";
            when "11" & x"57a" => DATA <= x"e706";
            when "11" & x"57b" => DATA <= x"0d00";
            when "11" & x"57c" => DATA <= x"07c0";
            when "11" & x"57d" => DATA <= x"e04a";
            when "11" & x"57e" => DATA <= x"0001";
            when "11" & x"57f" => DATA <= x"8008";
            when "11" & x"580" => DATA <= x"880e";
            when "11" & x"581" => DATA <= x"0008";
            when "11" & x"582" => DATA <= x"0010";
            when "11" & x"583" => DATA <= x"ef80";
            when "11" & x"584" => DATA <= x"0015";
            when "11" & x"585" => DATA <= x"83c0";
            when "11" & x"586" => DATA <= x"0072";
            when "11" & x"587" => DATA <= x"980c";
            when "11" & x"588" => DATA <= x"10c0";
            when "11" & x"589" => DATA <= x"e003";
            when "11" & x"58a" => DATA <= x"8008";
            when "11" & x"58b" => DATA <= x"0080";
            when "11" & x"58c" => DATA <= x"7fd0";
            when "11" & x"58d" => DATA <= x"013d";
            when "11" & x"58e" => DATA <= x"9e8f";
            when "11" & x"58f" => DATA <= x"0030";
            when "11" & x"590" => DATA <= x"5ff4";
            when "11" & x"591" => DATA <= x"0141";
            when "11" & x"592" => DATA <= x"23b0";
            when "11" & x"593" => DATA <= x"0381";
            when "11" & x"594" => DATA <= x"fec0";
            when "11" & x"595" => DATA <= x"2002";
            when "11" & x"596" => DATA <= x"000c";
            when "11" & x"597" => DATA <= x"8207";
            when "11" & x"598" => DATA <= x"0000";
            when "11" & x"599" => DATA <= x"c300";
            when "11" & x"59a" => DATA <= x"02ef";
            when "11" & x"59b" => DATA <= x"8000";
            when "11" & x"59c" => DATA <= x"6402";
            when "11" & x"59d" => DATA <= x"9802";
            when "11" & x"59e" => DATA <= x"0006";
            when "11" & x"59f" => DATA <= x"04c0";
            when "11" & x"5a0" => DATA <= x"7000";
            when "11" & x"5a1" => DATA <= x"1fc0";
            when "11" & x"5a2" => DATA <= x"3400";
            when "11" & x"5a3" => DATA <= x"0460";
            when "11" & x"5a4" => DATA <= x"a000";
            when "11" & x"5a5" => DATA <= x"8700";
            when "11" & x"5a6" => DATA <= x"0874";
            when "11" & x"5a7" => DATA <= x"0005";
            when "11" & x"5a8" => DATA <= x"4004";
            when "11" & x"5a9" => DATA <= x"f405";
            when "11" & x"5aa" => DATA <= x"8010";
            when "11" & x"5ab" => DATA <= x"3400";
            when "11" & x"5ac" => DATA <= x"05e0";
            when "11" & x"5ad" => DATA <= x"1200";
            when "11" & x"5ae" => DATA <= x"04a3";
            when "11" & x"5af" => DATA <= x"87c1";
            when "11" & x"5b0" => DATA <= x"82c0";
            when "11" & x"5b1" => DATA <= x"1fe5";
            when "11" & x"5b2" => DATA <= x"8d00";
            when "11" & x"5b3" => DATA <= x"083f";
            when "11" & x"5b4" => DATA <= x"dbfa";
            when "11" & x"5b5" => DATA <= x"0010";
            when "11" & x"5b6" => DATA <= x"7faf";
            when "11" & x"5b7" => DATA <= x"ec01";
            when "11" & x"5b8" => DATA <= x"fe10";
            when "11" & x"5b9" => DATA <= x"e080";
            when "11" & x"5ba" => DATA <= x"0570";
            when "11" & x"5bb" => DATA <= x"3ff4";
            when "11" & x"5bc" => DATA <= x"00be";
            when "11" & x"5bd" => DATA <= x"ac38";
            when "11" & x"5be" => DATA <= x"6803";
            when "11" & x"5bf" => DATA <= x"e063";
            when "11" & x"5c0" => DATA <= x"600e";
            when "11" & x"5c1" => DATA <= x"f575";
            when "11" & x"5c2" => DATA <= x"8000";
            when "11" & x"5c3" => DATA <= x"db76";
            when "11" & x"5c4" => DATA <= x"00cf";
            when "11" & x"5c5" => DATA <= x"0700";
            when "11" & x"5c6" => DATA <= x"1012";
            when "11" & x"5c7" => DATA <= x"0017";
            when "11" & x"5c8" => DATA <= x"0f00";
            when "11" & x"5c9" => DATA <= x"0040";
            when "11" & x"5ca" => DATA <= x"0025";
            when "11" & x"5cb" => DATA <= x"0001";
            when "11" & x"5cc" => DATA <= x"9880";
            when "11" & x"5cd" => DATA <= x"0008";
            when "11" & x"5ce" => DATA <= x"0007";
            when "11" & x"5cf" => DATA <= x"4004";
            when "11" & x"5d0" => DATA <= x"43e2";
            when "11" & x"5d1" => DATA <= x"5280";
            when "11" & x"5d2" => DATA <= x"020a";
            when "11" & x"5d3" => DATA <= x"9003";
            when "11" & x"5d4" => DATA <= x"05f6";
            when "11" & x"5d5" => DATA <= x"f2e0";
            when "11" & x"5d6" => DATA <= x"0008";
            when "11" & x"5d7" => DATA <= x"01c8";
            when "11" & x"5d8" => DATA <= x"ff53";
            when "11" & x"5d9" => DATA <= x"f003";
            when "11" & x"5da" => DATA <= x"0030";
            when "11" & x"5db" => DATA <= x"017f";
            when "11" & x"5dc" => DATA <= x"9958";
            when "11" & x"5dd" => DATA <= x"0100";
            when "11" & x"5de" => DATA <= x"f80e";
            when "11" & x"5df" => DATA <= x"801f";
            when "11" & x"5e0" => DATA <= x"e1f9";
            when "11" & x"5e1" => DATA <= x"0000";
            when "11" & x"5e2" => DATA <= x"b428";
            when "11" & x"5e3" => DATA <= x"01b9";
            when "11" & x"5e4" => DATA <= x"2000";
            when "11" & x"5e5" => DATA <= x"fa00";
            when "11" & x"5e6" => DATA <= x"6348";
            when "11" & x"5e7" => DATA <= x"0202";
            when "11" & x"5e8" => DATA <= x"8000";
            when "11" & x"5e9" => DATA <= x"8800";
            when "11" & x"5ea" => DATA <= x"002c";
            when "11" & x"5eb" => DATA <= x"01dc";
            when "11" & x"5ec" => DATA <= x"0804";
            when "11" & x"5ed" => DATA <= x"8341";
            when "11" & x"5ee" => DATA <= x"00d0";
            when "11" & x"5ef" => DATA <= x"aee2";
            when "11" & x"5f0" => DATA <= x"71ba";
            when "11" & x"5f1" => DATA <= x"938d";
            when "11" & x"5f2" => DATA <= x"e6e2";
            when "11" & x"5f3" => DATA <= x"bfaa";
            when "11" & x"5f4" => DATA <= x"dfab";
            when "11" & x"5f5" => DATA <= x"94ca";
            when "11" & x"5f6" => DATA <= x"caba";
            when "11" & x"5f7" => DATA <= x"a75a";
            when "11" & x"5f8" => DATA <= x"a914";
            when "11" & x"5f9" => DATA <= x"8041";
            when "11" & x"5fa" => DATA <= x"2a95";
            when "11" & x"5fb" => DATA <= x"6aa5";
            when "11" & x"5fc" => DATA <= x"5fbf";
            when "11" & x"5fd" => DATA <= x"9ff8";
            when "11" & x"5fe" => DATA <= x"018a";
            when "11" & x"5ff" => DATA <= x"c10c";
            when "11" & x"600" => DATA <= x"57c0";
            when "11" & x"601" => DATA <= x"11b0";
            when "11" & x"602" => DATA <= x"fc7f";
            when "11" & x"603" => DATA <= x"80c0";
            when "11" & x"604" => DATA <= x"0c77";
            when "11" & x"605" => DATA <= x"fa01";
            when "11" & x"606" => DATA <= x"0881";
            when "11" & x"607" => DATA <= x"4781";
            when "11" & x"608" => DATA <= x"c003";
            when "11" & x"609" => DATA <= x"fdff";
            when "11" & x"60a" => DATA <= x"7dd0";
            when "11" & x"60b" => DATA <= x"033f";
            when "11" & x"60c" => DATA <= x"7fda";
            when "11" & x"60d" => DATA <= x"0fb7";
            when "11" & x"60e" => DATA <= x"9f80";
            when "11" & x"60f" => DATA <= x"807c";
            when "11" & x"610" => DATA <= x"0000";
            when "11" & x"611" => DATA <= x"e076";
            when "11" & x"612" => DATA <= x"77fb";
            when "11" & x"613" => DATA <= x"bebf";
            when "11" & x"614" => DATA <= x"ecf9";
            when "11" & x"615" => DATA <= x"7e0f";
            when "11" & x"616" => DATA <= x"0008";
            when "11" & x"617" => DATA <= x"a802";
            when "11" & x"618" => DATA <= x"bf10";
            when "11" & x"619" => DATA <= x"3400";
            when "11" & x"61a" => DATA <= x"04a0";
            when "11" & x"61b" => DATA <= x"0aff";
            when "11" & x"61c" => DATA <= x"401e";
            when "11" & x"61d" => DATA <= x"1c0e";
            when "11" & x"61e" => DATA <= x"1603";
            when "11" & x"61f" => DATA <= x"b99e";
            when "11" & x"620" => DATA <= x"c773";
            when "11" & x"621" => DATA <= x"b838";
            when "11" & x"622" => DATA <= x"7d3e";
            when "11" & x"623" => DATA <= x"1f0d";
            when "11" & x"624" => DATA <= x"a7c3";
            when "11" & x"625" => DATA <= x"e052";
            when "11" & x"626" => DATA <= x"2904";
            when "11" & x"627" => DATA <= x"8000";
            when "11" & x"628" => DATA <= x"2211";
            when "11" & x"629" => DATA <= x"4892";
            when "11" & x"62a" => DATA <= x"fb3f";
            when "11" & x"62b" => DATA <= x"bda6";
            when "11" & x"62c" => DATA <= x"e573";
            when "11" & x"62d" => DATA <= x"3d8c";
            when "11" & x"62e" => DATA <= x"c7ea";
            when "11" & x"62f" => DATA <= x"0020";
            when "11" & x"630" => DATA <= x"adc9";
            when "11" & x"631" => DATA <= x"8ff0";
            when "11" & x"632" => DATA <= x"02ce";
            when "11" & x"633" => DATA <= x"8000";
            when "11" & x"634" => DATA <= x"4af1";
            when "11" & x"635" => DATA <= x"33fc";
            when "11" & x"636" => DATA <= x"00d9";
            when "11" & x"637" => DATA <= x"a004";
            when "11" & x"638" => DATA <= x"0b7d";
            when "11" & x"639" => DATA <= x"66ff";
            when "11" & x"63a" => DATA <= x"0033";
            when "11" & x"63b" => DATA <= x"3800";
            when "11" & x"63c" => DATA <= x"de99";
            when "11" & x"63d" => DATA <= x"7f80";
            when "11" & x"63e" => DATA <= x"04dc";
            when "11" & x"63f" => DATA <= x"00b3";
            when "11" & x"640" => DATA <= x"263f";
            when "11" & x"641" => DATA <= x"c00b";
            when "11" & x"642" => DATA <= x"3e00";
            when "11" & x"643" => DATA <= x"6a99";
            when "11" & x"644" => DATA <= x"9fe0";
            when "11" & x"645" => DATA <= x"04cf";
            when "11" & x"646" => DATA <= x"001e";
            when "11" & x"647" => DATA <= x"866f";
            when "11" & x"648" => DATA <= x"f003";
            when "11" & x"649" => DATA <= x"3400";
            when "11" & x"64a" => DATA <= x"6000";
            when "11" & x"64b" => DATA <= x"1b53";
            when "11" & x"64c" => DATA <= x"2ff0";
            when "11" & x"64d" => DATA <= x"0198";
            when "11" & x"64e" => DATA <= x"0004";
            when "11" & x"64f" => DATA <= x"1037";
            when "11" & x"650" => DATA <= x"8d8f";
            when "11" & x"651" => DATA <= x"f001";
            when "11" & x"652" => DATA <= x"be80";
            when "11" & x"653" => DATA <= x"0807";
            when "11" & x"654" => DATA <= x"f613";
            when "11" & x"655" => DATA <= x"fc00";
            when "11" & x"656" => DATA <= x"fe00";
            when "11" & x"657" => DATA <= x"3418";
            when "11" & x"658" => DATA <= x"0ef0";
            when "11" & x"659" => DATA <= x"b3fc";
            when "11" & x"65a" => DATA <= x"00b6";
            when "11" & x"65b" => DATA <= x"2850";
            when "11" & x"65c" => DATA <= x"03fd";
            when "11" & x"65d" => DATA <= x"f0ff";
            when "11" & x"65e" => DATA <= x"0024";
            when "11" & x"65f" => DATA <= x"4000";
            when "11" & x"660" => DATA <= x"8243";
            when "11" & x"661" => DATA <= x"fdde";
            when "11" & x"662" => DATA <= x"1d7c";
            when "11" & x"663" => DATA <= x"00c0";
            when "11" & x"664" => DATA <= x"0040";
            when "11" & x"665" => DATA <= x"3365";
            when "11" & x"666" => DATA <= x"fefe";
            when "11" & x"667" => DATA <= x"6f85";
            when "11" & x"668" => DATA <= x"4042";
            when "11" & x"669" => DATA <= x"0002";
            when "11" & x"66a" => DATA <= x"ffbf";
            when "11" & x"66b" => DATA <= x"f801";
            when "11" & x"66c" => DATA <= x"00f7";
            when "11" & x"66d" => DATA <= x"5fbf";
            when "11" & x"66e" => DATA <= x"d7f2";
            when "11" & x"66f" => DATA <= x"00fe";
            when "11" & x"670" => DATA <= x"7d8f";
            when "11" & x"671" => DATA <= x"dbe0";
            when "11" & x"672" => DATA <= x"07e0";
            when "11" & x"673" => DATA <= x"0c04";
            when "11" & x"674" => DATA <= x"ff7d";
            when "11" & x"675" => DATA <= x"bf03";
            when "11" & x"676" => DATA <= x"8001";
            when "11" & x"677" => DATA <= x"7811";
            when "11" & x"678" => DATA <= x"00d7";
            when "11" & x"679" => DATA <= x"7bb3";
            when "11" & x"67a" => DATA <= x"e800";
            when "11" & x"67b" => DATA <= x"04cc";
            when "11" & x"67c" => DATA <= x"003f";
            when "11" & x"67d" => DATA <= x"dfcf";
            when "11" & x"67e" => DATA <= x"b3e5";
            when "11" & x"67f" => DATA <= x"0004";
            when "11" & x"680" => DATA <= x"060f";
            when "11" & x"681" => DATA <= x"daff";
            when "11" & x"682" => DATA <= x"77d0";
            when "11" & x"683" => DATA <= x"0081";
            when "11" & x"684" => DATA <= x"467f";
            when "11" & x"685" => DATA <= x"7f83";
            when "11" & x"686" => DATA <= x"dff4";
            when "11" & x"687" => DATA <= x"00aa";
            when "11" & x"688" => DATA <= x"59d7";
            when "11" & x"689" => DATA <= x"f805";
            when "11" & x"68a" => DATA <= x"de00";
            when "11" & x"68b" => DATA <= x"782e";
            when "11" & x"68c" => DATA <= x"1166";
            when "11" & x"68d" => DATA <= x"b7f0";
            when "11" & x"68e" => DATA <= x"01ee";
            when "11" & x"68f" => DATA <= x"007f";
            when "11" & x"690" => DATA <= x"b058";
            when "11" & x"691" => DATA <= x"0fe7";
            when "11" & x"692" => DATA <= x"f801";
            when "11" & x"693" => DATA <= x"ea00";
            when "11" & x"694" => DATA <= x"7fb7";
            when "11" & x"695" => DATA <= x"0a0f";
            when "11" & x"696" => DATA <= x"f6f8";
            when "11" & x"697" => DATA <= x"01fe";
            when "11" & x"698" => DATA <= x"007f";
            when "11" & x"699" => DATA <= x"d003";
            when "11" & x"69a" => DATA <= x"fdfc";
            when "11" & x"69b" => DATA <= x"007f";
            when "11" & x"69c" => DATA <= x"8018";
            when "11" & x"69d" => DATA <= x"0011";
            when "11" & x"69e" => DATA <= x"057f";
            when "11" & x"69f" => DATA <= x"8017";
            when "11" & x"6a0" => DATA <= x"f400";
            when "11" & x"6a1" => DATA <= x"0200";
            when "11" & x"6a2" => DATA <= x"d7f8";
            when "11" & x"6a3" => DATA <= x"01fc";
            when "11" & x"6a4" => DATA <= x"40e0";
            when "11" & x"6a5" => DATA <= x"0aff";
            when "11" & x"6a6" => DATA <= x"003f";
            when "11" & x"6a7" => DATA <= x"f800";
            when "11" & x"6a8" => DATA <= x"415f";
            when "11" & x"6a9" => DATA <= x"e007";
            when "11" & x"6aa" => DATA <= x"ff00";
            when "11" & x"6ab" => DATA <= x"006b";
            when "11" & x"6ac" => DATA <= x"fc00";
            when "11" & x"6ad" => DATA <= x"ffe0";
            when "11" & x"6ae" => DATA <= x"0013";
            when "11" & x"6af" => DATA <= x"fd06";
            when "11" & x"6b0" => DATA <= x"005f";
            when "11" & x"6b1" => DATA <= x"d010";
            when "11" & x"6b2" => DATA <= x"00e0";
            when "11" & x"6b3" => DATA <= x"ff04";
            when "11" & x"6b4" => DATA <= x"a013";
            when "11" & x"6b5" => DATA <= x"e000";
            when "11" & x"6b6" => DATA <= x"6044";
            when "11" & x"6b7" => DATA <= x"8cff";
            when "11" & x"6b8" => DATA <= x"1980";
            when "11" & x"6b9" => DATA <= x"1f7c";
            when "11" & x"6ba" => DATA <= x"0050";
            when "11" & x"6bb" => DATA <= x"7f80";
            when "11" & x"6bc" => DATA <= x"080c";
            when "11" & x"6bd" => DATA <= x"fe00";
            when "11" & x"6be" => DATA <= x"0237";
            when "11" & x"6bf" => DATA <= x"c60f";
            when "11" & x"6c0" => DATA <= x"800b";
            when "11" & x"6c1" => DATA <= x"2380";
            when "11" & x"6c2" => DATA <= x"1d89";
            when "11" & x"6c3" => DATA <= x"97f8";
            when "11" & x"6c4" => DATA <= x"00c9";
            when "11" & x"6c5" => DATA <= x"4002";
            when "11" & x"6c6" => DATA <= x"03b3";
            when "11" & x"6c7" => DATA <= x"25fe";
            when "11" & x"6c8" => DATA <= x"0019";
            when "11" & x"6c9" => DATA <= x"5000";
            when "11" & x"6ca" => DATA <= x"8176";
            when "11" & x"6cb" => DATA <= x"647f";
            when "11" & x"6cc" => DATA <= x"8013";
            when "11" & x"6cd" => DATA <= x"6800";
            when "11" & x"6ce" => DATA <= x"0161";
            when "11" & x"6cf" => DATA <= x"fe56";
            when "11" & x"6d0" => DATA <= x"7fbc";
            when "11" & x"6d1" => DATA <= x"08b4";
            when "11" & x"6d2" => DATA <= x"00ad";
            when "11" & x"6d3" => DATA <= x"1ab2";
            when "11" & x"6d4" => DATA <= x"5bef";
            when "11" & x"6d5" => DATA <= x"f23d";
            when "11" & x"6d6" => DATA <= x"0001";
            when "11" & x"6d7" => DATA <= x"9fe8";
            when "11" & x"6d8" => DATA <= x"47fb";
            when "11" & x"6d9" => DATA <= x"3803";
            when "11" & x"6da" => DATA <= x"c00f";
            when "11" & x"6db" => DATA <= x"f093";
            when "11" & x"6dc" => DATA <= x"cd77";
            when "11" & x"6dd" => DATA <= x"c000";
            when "11" & x"6de" => DATA <= x"44a8";
            when "11" & x"6df" => DATA <= x"90fe";
            when "11" & x"6e0" => DATA <= x"fb00";
            when "11" & x"6e1" => DATA <= x"2400";
            when "11" & x"6e2" => DATA <= x"0807";
            when "11" & x"6e3" => DATA <= x"e822";
            when "11" & x"6e4" => DATA <= x"bfc0";
            when "11" & x"6e5" => DATA <= x"0420";
            when "11" & x"6e6" => DATA <= x"0045";
            when "11" & x"6e7" => DATA <= x"ee00";
            when "11" & x"6e8" => DATA <= x"7fbe";
            when "11" & x"6e9" => DATA <= x"4000";
            when "11" & x"6ea" => DATA <= x"8000";
            when "11" & x"6eb" => DATA <= x"99fe";
            when "11" & x"6ec" => DATA <= x"067f";
            when "11" & x"6ed" => DATA <= x"bbe4";
            when "11" & x"6ee" => DATA <= x"01fe";
            when "11" & x"6ef" => DATA <= x"247f";
            when "11" & x"6f0" => DATA <= x"bf38";
            when "11" & x"6f1" => DATA <= x"0100";
            when "11" & x"6f2" => DATA <= x"ff50";
            when "11" & x"6f3" => DATA <= x"57ff";
            when "11" & x"6f4" => DATA <= x"000e";
            when "11" & x"6f5" => DATA <= x"1fe0";
            when "11" & x"6f6" => DATA <= x"0aff";
            when "11" & x"6f7" => DATA <= x"0000";
            when "11" & x"6f8" => DATA <= x"8002";
            when "11" & x"6f9" => DATA <= x"0338";
            when "11" & x"6fa" => DATA <= x"01ec";
            when "11" & x"6fb" => DATA <= x"7690";
            when "11" & x"6fc" => DATA <= x"07f9";
            when "11" & x"6fd" => DATA <= x"41fe";
            when "11" & x"6fe" => DATA <= x"7fe0";
            when "11" & x"6ff" => DATA <= x"0061";
            when "11" & x"700" => DATA <= x"fc08";
            when "11" & x"701" => DATA <= x"7f77";
            when "11" & x"702" => DATA <= x"c803";
            when "11" & x"703" => DATA <= x"dc00";
            when "11" & x"704" => DATA <= x"fb5b";
            when "11" & x"705" => DATA <= x"c803";
            when "11" & x"706" => DATA <= x"6c44";
            when "11" & x"707" => DATA <= x"f77f";
            when "11" & x"708" => DATA <= x"f003";
            when "11" & x"709" => DATA <= x"91fe";
            when "11" & x"70a" => DATA <= x"007f";
            when "11" & x"70b" => DATA <= x"ae40";
            when "11" & x"70c" => DATA <= x"14e0";
            when "11" & x"70d" => DATA <= x"7e3e";
            when "11" & x"70e" => DATA <= x"802b";
            when "11" & x"70f" => DATA <= x"fde0";
            when "11" & x"710" => DATA <= x"0f37";
            when "11" & x"711" => DATA <= x"93cd";
            when "11" & x"712" => DATA <= x"eef0";
            when "11" & x"713" => DATA <= x"fbfc";
            when "11" & x"714" => DATA <= x"7e55";
            when "11" & x"715" => DATA <= x"2a72";
            when "11" & x"716" => DATA <= x"a800";
            when "11" & x"717" => DATA <= x"ae00";
            when "11" & x"718" => DATA <= x"3ab9";
            when "11" & x"719" => DATA <= x"4ca7";
            when "11" & x"71a" => DATA <= x"57aa";
            when "11" & x"71b" => DATA <= x"c15e";
            when "11" & x"71c" => DATA <= x"0045";
            when "11" & x"71d" => DATA <= x"0294";
            when "11" & x"71e" => DATA <= x"0f05";
            when "11" & x"71f" => DATA <= x"331c";
            when "11" & x"720" => DATA <= x"4f55";
            when "11" & x"721" => DATA <= x"eb05";
            when "11" & x"722" => DATA <= x"6a2d";
            when "11" & x"723" => DATA <= x"56af";
            when "11" & x"724" => DATA <= x"7f3a";
            when "11" & x"725" => DATA <= x"48f4";
            when "11" & x"726" => DATA <= x"feff";
            when "11" & x"727" => DATA <= x"a7f6";
            when "11" & x"728" => DATA <= x"39fc";
            when "11" & x"729" => DATA <= x"0010";
            when "11" & x"72a" => DATA <= x"003e";
            when "11" & x"72b" => DATA <= x"c000";
            when "11" & x"72c" => DATA <= x"8013";
            when "11" & x"72d" => DATA <= x"e380";
            when "11" & x"72e" => DATA <= x"007c";
            when "11" & x"72f" => DATA <= x"00ff";
            when "11" & x"730" => DATA <= x"7000";
            when "11" & x"731" => DATA <= x"2a02";
            when "11" & x"732" => DATA <= x"801c";
            when "11" & x"733" => DATA <= x"1fff";
            when "11" & x"734" => DATA <= x"5ff5";
            when "11" & x"735" => DATA <= x"f77f";
            when "11" & x"736" => DATA <= x"fe02";
            when "11" & x"737" => DATA <= x"01f0";
            when "11" & x"738" => DATA <= x"0001";
            when "11" & x"739" => DATA <= x"bc0e";
            when "11" & x"73a" => DATA <= x"e103";
            when "11" & x"73b" => DATA <= x"b85d";
            when "11" & x"73c" => DATA <= x"8ef7";
            when "11" & x"73d" => DATA <= x"f801";
            when "11" & x"73e" => DATA <= x"00a0";
            when "11" & x"73f" => DATA <= x"5e0f";
            when "11" & x"740" => DATA <= x"baf9";
            when "11" & x"741" => DATA <= x"fd60";
            when "11" & x"742" => DATA <= x"15ff";
            when "11" & x"743" => DATA <= x"600f";
            when "11" & x"744" => DATA <= x"f603";
            when "11" & x"745" => DATA <= x"8001";
            when "11" & x"746" => DATA <= x"5c4c";
            when "11" & x"747" => DATA <= x"2703";
            when "11" & x"748" => DATA <= x"003d";
            when "11" & x"749" => DATA <= x"c3e9";
            when "11" & x"74a" => DATA <= x"fa1f";
            when "11" & x"74b" => DATA <= x"0f11";
            when "11" & x"74c" => DATA <= x"081c";
            when "11" & x"74d" => DATA <= x"8a05";
            when "11" & x"74e" => DATA <= x"2215";
            when "11" & x"74f" => DATA <= x"abf6";
            when "11" & x"750" => DATA <= x"8078";
            when "11" & x"751" => DATA <= x"0080";
            when "11" & x"752" => DATA <= x"007f";
            when "11" & x"753" => DATA <= x"bf8f";
            when "11" & x"754" => DATA <= x"d3fc";
            when "11" & x"755" => DATA <= x"2d5d";
            when "11" & x"756" => DATA <= x"c802";
            when "11" & x"757" => DATA <= x"e000";
            when "11" & x"758" => DATA <= x"eb6c";
            when "11" & x"759" => DATA <= x"c803";
            when "11" & x"75a" => DATA <= x"7400";
            when "11" & x"75b" => DATA <= x"5876";
            when "11" & x"75c" => DATA <= x"4803";
            when "11" & x"75d" => DATA <= x"bc00";
            when "11" & x"75e" => DATA <= x"a933";
            when "11" & x"75f" => DATA <= x"4801";
            when "11" & x"760" => DATA <= x"f800";
            when "11" & x"761" => DATA <= x"da5b";
            when "11" & x"762" => DATA <= x"c802";
            when "11" & x"763" => DATA <= x"fc00";
            when "11" & x"764" => DATA <= x"bd4c";
            when "11" & x"765" => DATA <= x"c803";
            when "11" & x"766" => DATA <= x"7c00";
            when "11" & x"767" => DATA <= x"7f66";
            when "11" & x"768" => DATA <= x"c803";
            when "11" & x"769" => DATA <= x"f400";
            when "11" & x"76a" => DATA <= x"bd33";
            when "11" & x"76b" => DATA <= x"4801";
            when "11" & x"76c" => DATA <= x"1800";
            when "11" & x"76d" => DATA <= x"563f";
            when "11" & x"76e" => DATA <= x"c800";
            when "11" & x"76f" => DATA <= x"4400";
            when "11" & x"770" => DATA <= x"6776";
            when "11" & x"771" => DATA <= x"5800";
            when "11" & x"772" => DATA <= x"7477";
            when "11" & x"773" => DATA <= x"6008";
            when "11" & x"774" => DATA <= x"0678";
            when "11" & x"775" => DATA <= x"8280";
            when "11" & x"776" => DATA <= x"0400";
            when "11" & x"777" => DATA <= x"0080";
            when "11" & x"778" => DATA <= x"1059";
            when "11" & x"779" => DATA <= x"e00f";
            when "11" & x"77a" => DATA <= x"f000";
            when "11" & x"77b" => DATA <= x"4240";
            when "11" & x"77c" => DATA <= x"092f";
            when "11" & x"77d" => DATA <= x"f000";
            when "11" & x"77e" => DATA <= x"8240";
            when "11" & x"77f" => DATA <= x"0681";
            when "11" & x"780" => DATA <= x"c000";
            when "11" & x"781" => DATA <= x"5680";
            when "11" & x"782" => DATA <= x"0600";
            when "11" & x"783" => DATA <= x"0022";
            when "11" & x"784" => DATA <= x"0400";
            when "11" & x"785" => DATA <= x"20a0";
            when "11" & x"786" => DATA <= x"0510";
            when "11" & x"787" => DATA <= x"0806";
            when "11" & x"788" => DATA <= x"dbb0";
            when "11" & x"789" => DATA <= x"0021";
            when "11" & x"78a" => DATA <= x"d440";
            when "11" & x"78b" => DATA <= x"4001";
            when "11" & x"78c" => DATA <= x"0808";
            when "11" & x"78d" => DATA <= x"0030";
            when "11" & x"78e" => DATA <= x"e3aa";
            when "11" & x"78f" => DATA <= x"80a8";
            when "11" & x"790" => DATA <= x"0004";
            when "11" & x"791" => DATA <= x"0017";
            when "11" & x"792" => DATA <= x"16c4";
            when "11" & x"793" => DATA <= x"5600";
            when "11" & x"794" => DATA <= x"6fb0";
            when "11" & x"795" => DATA <= x"0403";
            when "11" & x"796" => DATA <= x"7f40";
            when "11" & x"797" => DATA <= x"0020";
            when "11" & x"798" => DATA <= x"37e2";
            when "11" & x"799" => DATA <= x"0240";
            when "11" & x"79a" => DATA <= x"0422";
            when "11" & x"79b" => DATA <= x"0338";
            when "11" & x"79c" => DATA <= x"0d00";
            when "11" & x"79d" => DATA <= x"0000";
            when "11" & x"79e" => DATA <= x"a000";
            when "11" & x"79f" => DATA <= x"0166";
            when "11" & x"7a0" => DATA <= x"3f80";
            when "11" & x"7a1" => DATA <= x"28e4";
            when "11" & x"7a2" => DATA <= x"01e4";
            when "11" & x"7a3" => DATA <= x"0040";
            when "11" & x"7a4" => DATA <= x"1fa4";
            when "11" & x"7a5" => DATA <= x"00fe";
            when "11" & x"7a6" => DATA <= x"0036";
            when "11" & x"7a7" => DATA <= x"0ce4";
            when "11" & x"7a8" => DATA <= x"017e";
            when "11" & x"7a9" => DATA <= x"0057";
            when "11" & x"7aa" => DATA <= x"b664";
            when "11" & x"7ab" => DATA <= x"01fe";
            when "11" & x"7ac" => DATA <= x"002d";
            when "11" & x"7ad" => DATA <= x"3364";
            when "11" & x"7ae" => DATA <= x"01fa";
            when "11" & x"7af" => DATA <= x"0052";
            when "11" & x"7b0" => DATA <= x"99a4";
            when "11" & x"7b1" => DATA <= x"007c";
            when "11" & x"7b2" => DATA <= x"0003";
            when "11" & x"7b3" => DATA <= x"3efc";
            when "11" & x"7b4" => DATA <= x"01f7";
            when "11" & x"7b5" => DATA <= x"200a";
            when "11" & x"7b6" => DATA <= x"0a00";
            when "11" & x"7b7" => DATA <= x"2980";
            when "11" & x"7b8" => DATA <= x"0214";
            when "11" & x"7b9" => DATA <= x"0010";
            when "11" & x"7ba" => DATA <= x"0008";
            when "11" & x"7bb" => DATA <= x"0ec0";
            when "11" & x"7bc" => DATA <= x"000c";
            when "11" & x"7bd" => DATA <= x"8014";
            when "11" & x"7be" => DATA <= x"19f2";
            when "11" & x"7bf" => DATA <= x"0084";
            when "11" & x"7c0" => DATA <= x"0021";
            when "11" & x"7c1" => DATA <= x"4c92";
            when "11" & x"7c2" => DATA <= x"006e";
            when "11" & x"7c3" => DATA <= x"0012";
            when "11" & x"7c4" => DATA <= x"86f2";
            when "11" & x"7c5" => DATA <= x"00f7";
            when "11" & x"7c6" => DATA <= x"0025";
            when "11" & x"7c7" => DATA <= x"5372";
            when "11" & x"7c8" => DATA <= x"00fb";
            when "11" & x"7c9" => DATA <= x"001e";
            when "11" & x"7ca" => DATA <= x"8fb4";
            when "11" & x"7cb" => DATA <= x"0080";
            when "11" & x"7cc" => DATA <= x"0001";
            when "11" & x"7cd" => DATA <= x"400f";
            when "11" & x"7ce" => DATA <= x"c3ed";
            when "11" & x"7cf" => DATA <= x"0600";
            when "11" & x"7d0" => DATA <= x"4294";
            when "11" & x"7d1" => DATA <= x"0850";
            when "11" & x"7d2" => DATA <= x"42d0";
            when "11" & x"7d3" => DATA <= x"0013";
            when "11" & x"7d4" => DATA <= x"8019";
            when "11" & x"7d5" => DATA <= x"0fd0";
            when "11" & x"7d6" => DATA <= x"00f0";
            when "11" & x"7d7" => DATA <= x"0014";
            when "11" & x"7d8" => DATA <= x"120f";
            when "11" & x"7d9" => DATA <= x"022f";
            when "11" & x"7da" => DATA <= x"bb00";
            when "11" & x"7db" => DATA <= x"6837";
            when "11" & x"7dc" => DATA <= x"821c";
            when "11" & x"7dd" => DATA <= x"0010";
            when "11" & x"7de" => DATA <= x"002e";
            when "11" & x"7df" => DATA <= x"5bf2";
            when "11" & x"7e0" => DATA <= x"0008";
            when "11" & x"7e1" => DATA <= x"000c";
            when "11" & x"7e2" => DATA <= x"59cc";
            when "11" & x"7e3" => DATA <= x"00c0";
            when "11" & x"7e4" => DATA <= x"0101";
            when "11" & x"7e5" => DATA <= x"4000";
            when "11" & x"7e6" => DATA <= x"14b5";
            when "11" & x"7e7" => DATA <= x"800c";
            when "11" & x"7e8" => DATA <= x"00fc";
            when "11" & x"7e9" => DATA <= x"0080";
            when "11" & x"7ea" => DATA <= x"a006";
            when "11" & x"7eb" => DATA <= x"3b00";
            when "11" & x"7ec" => DATA <= x"0340";
            when "11" & x"7ed" => DATA <= x"020a";
            when "11" & x"7ee" => DATA <= x"0020";
            when "11" & x"7ef" => DATA <= x"6800";
            when "11" & x"7f0" => DATA <= x"6000";
            when "11" & x"7f1" => DATA <= x"46a0";
            when "11" & x"7f2" => DATA <= x"010c";
            when "11" & x"7f3" => DATA <= x"8011";
            when "11" & x"7f4" => DATA <= x"1e60";
            when "11" & x"7f5" => DATA <= x"8008";
            when "11" & x"7f6" => DATA <= x"0011";
            when "11" & x"7f7" => DATA <= x"400c";
            when "11" & x"7f8" => DATA <= x"05f8";
            when "11" & x"7f9" => DATA <= x"103c";
            when "11" & x"7fa" => DATA <= x"0006";
            when "11" & x"7fb" => DATA <= x"0780";
            when "11" & x"7fc" => DATA <= x"02b1";
            when "11" & x"7fd" => DATA <= x"7780";
            when "11" & x"7fe" => DATA <= x"0216";
            when "11" & x"7ff" => DATA <= x"0080";
            when "11" & x"800" => DATA <= x"0282";
            when "11" & x"801" => DATA <= x"802b";
            when "11" & x"802" => DATA <= x"c1fc";
            when "11" & x"803" => DATA <= x"e8af";
            when "11" & x"804" => DATA <= x"8773";
            when "11" & x"805" => DATA <= x"f17f";
            when "11" & x"806" => DATA <= x"e7e0";
            when "11" & x"807" => DATA <= x"e3f0";
            when "11" & x"808" => DATA <= x"0168";
            when "11" & x"809" => DATA <= x"ff00";
            when "11" & x"80a" => DATA <= x"57fb";
            when "11" & x"80b" => DATA <= x"81e8";
            when "11" & x"80c" => DATA <= x"10ae";
            when "11" & x"80d" => DATA <= x"b005";
            when "11" & x"80e" => DATA <= x"55af";
            when "11" & x"80f" => DATA <= x"15ca";
            when "11" & x"810" => DATA <= x"8670";
            when "11" & x"811" => DATA <= x"b950";
            when "11" & x"812" => DATA <= x"b244";
            when "11" & x"813" => DATA <= x"3a55";
            when "11" & x"814" => DATA <= x"0aa4";
            when "11" & x"815" => DATA <= x"1201";
            when "11" & x"816" => DATA <= x"c551";
            when "11" & x"817" => DATA <= x"54fe";
            when "11" & x"818" => DATA <= x"3fd7";
            when "11" & x"819" => DATA <= x"fa08";
            when "11" & x"81a" => DATA <= x"60b1";
            when "11" & x"81b" => DATA <= x"6800";
            when "11" & x"81c" => DATA <= x"05c0";
            when "11" & x"81d" => DATA <= x"15fe";
            when "11" & x"81e" => DATA <= x"fc00";
            when "11" & x"81f" => DATA <= x"0100";
            when "11" & x"820" => DATA <= x"03e0";
            when "11" & x"821" => DATA <= x"001d";
            when "11" & x"822" => DATA <= x"1e81";
            when "11" & x"823" => DATA <= x"a800";
            when "11" & x"824" => DATA <= x"03bd";
            when "11" & x"825" => DATA <= x"00c0";
            when "11" & x"826" => DATA <= x"65bb";
            when "11" & x"827" => DATA <= x"fbfd";
            when "11" & x"828" => DATA <= x"f6f3";
            when "11" & x"829" => DATA <= x"69d7";
            when "11" & x"82a" => DATA <= x"9d7d";
            when "11" & x"82b" => DATA <= x"bffc";
            when "11" & x"82c" => DATA <= x"0403";
            when "11" & x"82d" => DATA <= x"4001";
            when "11" & x"82e" => DATA <= x"8d00";
            when "11" & x"82f" => DATA <= x"eff1";
            when "11" & x"830" => DATA <= x"7a1c";
            when "11" & x"831" => DATA <= x"db5c";
            when "11" & x"832" => DATA <= x"ebe5";
            when "11" & x"833" => DATA <= x"f81f";
            when "11" & x"834" => DATA <= x"8007";
            when "11" & x"835" => DATA <= x"83e3";
            when "11" & x"836" => DATA <= x"f80c";
            when "11" & x"837" => DATA <= x"00fc";
            when "11" & x"838" => DATA <= x"900a";
            when "11" & x"839" => DATA <= x"c07f";
            when "11" & x"83a" => DATA <= x"3fe4";
            when "11" & x"83b" => DATA <= x"01c0";
            when "11" & x"83c" => DATA <= x"e373";
            when "11" & x"83d" => DATA <= x"b3dc";
            when "11" & x"83e" => DATA <= x"c02a";
            when "11" & x"83f" => DATA <= x"e00b";
            when "11" & x"840" => DATA <= x"a7c3";
            when "11" & x"841" => DATA <= x"61f4";
            when "11" & x"842" => DATA <= x"f83e";
            when "11" & x"843" => DATA <= x"a7f9";
            when "11" & x"844" => DATA <= x"54a8";
            when "11" & x"845" => DATA <= x"56e5";
            when "11" & x"846" => DATA <= x"5a00";
            when "11" & x"847" => DATA <= x"2018";
            when "11" & x"848" => DATA <= x"0900";
            when "11" & x"849" => DATA <= x"0381";
            when "11" & x"84a" => DATA <= x"537f";
            when "11" & x"84b" => DATA <= x"8fd5";
            when "11" & x"84c" => DATA <= x"fdc0";
            when "11" & x"84d" => DATA <= x"001a";
            when "11" & x"84e" => DATA <= x"0008";
            when "11" & x"84f" => DATA <= x"4802";
            when "11" & x"850" => DATA <= x"0680";
            when "11" & x"851" => DATA <= x"0114";
            when "11" & x"852" => DATA <= x"00a1";
            when "11" & x"853" => DATA <= x"0010";
            when "11" & x"854" => DATA <= x"2800";
            when "11" & x"855" => DATA <= x"0940";
            when "11" & x"856" => DATA <= x"0d00";
            when "11" & x"857" => DATA <= x"0082";
            when "11" & x"858" => DATA <= x"8000";
            when "11" & x"859" => DATA <= x"9400";
            when "11" & x"85a" => DATA <= x"6800";
            when "11" & x"85b" => DATA <= x"0428";
            when "11" & x"85c" => DATA <= x"0005";
            when "11" & x"85d" => DATA <= x"4002";
            when "11" & x"85e" => DATA <= x"c000";
            when "11" & x"85f" => DATA <= x"2280";
            when "11" & x"860" => DATA <= x"1034";
            when "11" & x"861" => DATA <= x"0002";
            when "11" & x"862" => DATA <= x"0002";
            when "11" & x"863" => DATA <= x"2800";
            when "11" & x"864" => DATA <= x"8140";
            when "11" & x"865" => DATA <= x"00a0";
            when "11" & x"866" => DATA <= x"0012";
            when "11" & x"867" => DATA <= x"8004";
            when "11" & x"868" => DATA <= x"1400";
            when "11" & x"869" => DATA <= x"1000";
            when "11" & x"86a" => DATA <= x"00bc";
            when "11" & x"86b" => DATA <= x"0000";
            when "11" & x"86c" => DATA <= x"20b0";
            when "11" & x"86d" => DATA <= x"0015";
            when "11" & x"86e" => DATA <= x"0000";
            when "11" & x"86f" => DATA <= x"8000";
            when "11" & x"870" => DATA <= x"2a00";
            when "11" & x"871" => DATA <= x"0970";
            when "11" & x"872" => DATA <= x"0083";
            when "11" & x"873" => DATA <= x"8018";
            when "11" & x"874" => DATA <= x"1400";
            when "11" & x"875" => DATA <= x"4490";
            when "11" & x"876" => DATA <= x"0087";
            when "11" & x"877" => DATA <= x"8020";
            when "11" & x"878" => DATA <= x"3400";
            when "11" & x"879" => DATA <= x"2000";
            when "11" & x"87a" => DATA <= x"0248";
            when "11" & x"87b" => DATA <= x"0088";
            when "11" & x"87c" => DATA <= x"0002";
            when "11" & x"87d" => DATA <= x"1150";
            when "11" & x"87e" => DATA <= x"0202";
            when "11" & x"87f" => DATA <= x"4002";
            when "11" & x"880" => DATA <= x"1400";
            when "11" & x"881" => DATA <= x"18a0";
            when "11" & x"882" => DATA <= x"0100";
            when "11" & x"883" => DATA <= x"0005";
            when "11" & x"884" => DATA <= x"4000";
            when "11" & x"885" => DATA <= x"1580";
            when "11" & x"886" => DATA <= x"0005";
            when "11" & x"887" => DATA <= x"c000";
            when "11" & x"888" => DATA <= x"2f00";
            when "11" & x"889" => DATA <= x"0000";
            when "11" & x"88a" => DATA <= x"bc00";
            when "11" & x"88b" => DATA <= x"0520";
            when "11" & x"88c" => DATA <= x"008a";
            when "11" & x"88d" => DATA <= x"0040";
            when "11" & x"88e" => DATA <= x"7000";
            when "11" & x"88f" => DATA <= x"8c07";
            when "11" & x"890" => DATA <= x"e008";
            when "11" & x"891" => DATA <= x"a040";
            when "11" & x"892" => DATA <= x"01c4";
            when "11" & x"893" => DATA <= x"23e0";
            when "11" & x"894" => DATA <= x"0205";
            when "11" & x"895" => DATA <= x"8001";
            when "11" & x"896" => DATA <= x"3c02";
            when "11" & x"897" => DATA <= x"4004";
            when "11" & x"898" => DATA <= x"1400";
            when "11" & x"899" => DATA <= x"8490";
            when "11" & x"89a" => DATA <= x"0085";
            when "11" & x"89b" => DATA <= x"0010";
            when "11" & x"89c" => DATA <= x"8008";
            when "11" & x"89d" => DATA <= x"1a00";
            when "11" & x"89e" => DATA <= x"0450";
            when "11" & x"89f" => DATA <= x"02cc";
            when "11" & x"8a0" => DATA <= x"0040";
            when "11" & x"8a1" => DATA <= x"d000";
            when "11" & x"8a2" => DATA <= x"0800";
            when "11" & x"8a3" => DATA <= x"4140";
            when "11" & x"8a4" => DATA <= x"0049";
            when "11" & x"8a5" => DATA <= x"0012";
            when "11" & x"8a6" => DATA <= x"5000";
            when "11" & x"8a7" => DATA <= x"8240";
            when "11" & x"8a8" => DATA <= x"003a";
            when "11" & x"8a9" => DATA <= x"0010";
            when "11" & x"8aa" => DATA <= x"f00a";
            when "11" & x"8ab" => DATA <= x"0001";
            when "11" & x"8ac" => DATA <= x"6802";
            when "11" & x"8ad" => DATA <= x"0000";
            when "11" & x"8ae" => DATA <= x"40d0";
            when "11" & x"8af" => DATA <= x"058c";
            when "11" & x"8b0" => DATA <= x"8001";
            when "11" & x"8b1" => DATA <= x"2800";
            when "11" & x"8b2" => DATA <= x"b200";
            when "11" & x"8b3" => DATA <= x"1050";
            when "11" & x"8b4" => DATA <= x"000a";
            when "11" & x"8b5" => DATA <= x"8009";
            when "11" & x"8b6" => DATA <= x"8000";
            when "11" & x"8b7" => DATA <= x"8500";
            when "11" & x"8b8" => DATA <= x"2068";
            when "11" & x"8b9" => DATA <= x"0009";
            when "11" & x"8ba" => DATA <= x"4112";
            when "11" & x"8bb" => DATA <= x"0001";
            when "11" & x"8bc" => DATA <= x"d000";
            when "11" & x"8bd" => DATA <= x"0f80";
            when "11" & x"8be" => DATA <= x"0100";
            when "11" & x"8bf" => DATA <= x"0080";
            when "11" & x"8c0" => DATA <= x"80e0";
            when "11" & x"8c1" => DATA <= x"0020";
            when "11" & x"8c2" => DATA <= x"a003";
            when "11" & x"8c3" => DATA <= x"8700";
            when "11" & x"8c4" => DATA <= x"10a8";
            when "11" & x"8c5" => DATA <= x"0084";
            when "11" & x"8c6" => DATA <= x"0040";
            when "11" & x"8c7" => DATA <= x"0004";
            when "11" & x"8c8" => DATA <= x"040e";
            when "11" & x"8c9" => DATA <= x"0008";
            when "11" & x"8ca" => DATA <= x"7800";
            when "11" & x"8cb" => DATA <= x"4380";
            when "11" & x"8cc" => DATA <= x"1894";
            when "11" & x"8cd" => DATA <= x"0080";
            when "11" & x"8ce" => DATA <= x"6078";
            when "11" & x"8cf" => DATA <= x"0700";
            when "11" & x"8d0" => DATA <= x"1001";
            when "11" & x"8d1" => DATA <= x"5c00";
            when "11" & x"8d2" => DATA <= x"01e0";
            when "11" & x"8d3" => DATA <= x"041f";
            when "11" & x"8d4" => DATA <= x"0000";
            when "11" & x"8d5" => DATA <= x"7c01";
            when "11" & x"8d6" => DATA <= x"4140";
            when "11" & x"8d7" => DATA <= x"0203";
            when "11" & x"8d8" => DATA <= x"0000";
            when "11" & x"8d9" => DATA <= x"0340";
            when "11" & x"8da" => DATA <= x"0080";
            when "11" & x"8db" => DATA <= x"0004";
            when "11" & x"8dc" => DATA <= x"4000";
            when "11" & x"8dd" => DATA <= x"0080";
            when "11" & x"8de" => DATA <= x"011c";
            when "11" & x"8df" => DATA <= x"001e";
            when "11" & x"8e0" => DATA <= x"0050";
            when "11" & x"8e1" => DATA <= x"7012";
            when "11" & x"8e2" => DATA <= x"c001";
            when "11" & x"8e3" => DATA <= x"1200";
            when "11" & x"8e4" => DATA <= x"28a0";
            when "11" & x"8e5" => DATA <= x"8145";
            when "11" & x"8e6" => DATA <= x"7c3f";
            when "11" & x"8e7" => DATA <= x"abe1";
            when "11" & x"8e8" => DATA <= x"fce8";
            when "11" & x"8e9" => DATA <= x"7c3f";
            when "11" & x"8ea" => DATA <= x"f4fd";
            when "11" & x"8eb" => DATA <= x"7f47";
            when "11" & x"8ec" => DATA <= x"e00a";
            when "11" & x"8ed" => DATA <= x"ff00";
            when "11" & x"8ee" => DATA <= x"3feb";
            when "11" & x"8ef" => DATA <= x"fa80";
            when "11" & x"8f0" => DATA <= x"01ee";
            when "11" & x"8f1" => DATA <= x"f601";
            when "11" & x"8f2" => DATA <= x"2cde";
            when "11" & x"8f3" => DATA <= x"6b00";
            when "11" & x"8f4" => DATA <= x"5141";
            when "11" & x"8f5" => DATA <= x"228a";
            when "11" & x"8f6" => DATA <= x"05e0";
            when "11" & x"8f7" => DATA <= x"000a";
            when "11" & x"8f8" => DATA <= x"2aaa";
            when "11" & x"8f9" => DATA <= x"aa05";
            when "11" & x"8fa" => DATA <= x"54a3";
            when "11" & x"8fb" => DATA <= x"547b";
            when "11" & x"8fc" => DATA <= x"f9fc";
            when "11" & x"8fd" => DATA <= x"41c0";
            when "11" & x"8fe" => DATA <= x"0c50";
            when "11" & x"8ff" => DATA <= x"0861";
            when "11" & x"900" => DATA <= x"f000";
            when "11" & x"901" => DATA <= x"0212";
            when "11" & x"902" => DATA <= x"1f8f";
            when "11" & x"903" => DATA <= x"f400";
            when "11" & x"904" => DATA <= x"000f";
            when "11" & x"905" => DATA <= x"d008";
            when "11" & x"906" => DATA <= x"1a8f";
            when "11" & x"907" => DATA <= x"a00b";
            when "11" & x"908" => DATA <= x"ff64";
            when "11" & x"909" => DATA <= x"002f";
            when "11" & x"90a" => DATA <= x"fdf6";
            when "11" & x"90b" => DATA <= x"f300";
            when "11" & x"90c" => DATA <= x"eb8d";
            when "11" & x"90d" => DATA <= x"00e8";
            when "11" & x"90e" => DATA <= x"0508";
            when "11" & x"90f" => DATA <= x"003b";
            when "11" & x"910" => DATA <= x"bfbf";
            when "11" & x"911" => DATA <= x"dde2";
            when "11" & x"912" => DATA <= x"793e";
            when "11" & x"913" => DATA <= x"5f8f";
            when "11" & x"914" => DATA <= x"e402";
            when "11" & x"915" => DATA <= x"bf00";
            when "11" & x"916" => DATA <= x"e007";
            when "11" & x"917" => DATA <= x"8700";
            when "11" & x"918" => DATA <= x"3fd9";
            when "11" & x"919" => DATA <= x"ec03";
            when "11" & x"91a" => DATA <= x"e3fc";
            when "11" & x"91b" => DATA <= x"0080";
            when "11" & x"91c" => DATA <= x"7332";
            when "11" & x"91d" => DATA <= x"d8ee";
            when "11" & x"91e" => DATA <= x"7703";
            when "11" & x"91f" => DATA <= x"01c0";
            when "11" & x"920" => DATA <= x"1f4f";
            when "11" & x"921" => DATA <= x"87c3";
            when "11" & x"922" => DATA <= x"69f0";
            when "11" & x"923" => DATA <= x"b878";
            when "11" & x"924" => DATA <= x"3e51";
            when "11" & x"925" => DATA <= x"2914";
            when "11" & x"926" => DATA <= x"0281";
            when "11" & x"927" => DATA <= x"5a14";
            when "11" & x"928" => DATA <= x"a002";
            when "11" & x"929" => DATA <= x"8500";
            when "11" & x"92a" => DATA <= x"1528";
            when "11" & x"92b" => DATA <= x"00a9";
            when "11" & x"92c" => DATA <= x"ffcf";
            when "11" & x"92d" => DATA <= x"ee00";
            when "11" & x"92e" => DATA <= x"5c78";
            when "11" & x"92f" => DATA <= x"037f";
            when "11" & x"930" => DATA <= x"c01f";
            when "11" & x"931" => DATA <= x"fe00";
            when "11" & x"932" => DATA <= x"7fa0";
            when "11" & x"933" => DATA <= x"0084";
            when "11" & x"934" => DATA <= x"802f";
            when "11" & x"935" => DATA <= x"e800";
            when "11" & x"936" => DATA <= x"1120";
            when "11" & x"937" => DATA <= x"0dff";
            when "11" & x"938" => DATA <= x"007e";
            when "11" & x"939" => DATA <= x"f803";
            when "11" & x"93a" => DATA <= x"fbc0";
            when "11" & x"93b" => DATA <= x"0234";
            when "11" & x"93c" => DATA <= x"0010";
            when "11" & x"93d" => DATA <= x"f00f";
            when "11" & x"93e" => DATA <= x"00d0";
            when "11" & x"93f" => DATA <= x"0010";
            when "11" & x"940" => DATA <= x"0020";
            when "11" & x"941" => DATA <= x"0210";
            when "11" & x"942" => DATA <= x"7002";
            when "11" & x"943" => DATA <= x"03c0";
            when "11" & x"944" => DATA <= x"3c03";
            when "11" & x"945" => DATA <= x"c002";
            when "11" & x"946" => DATA <= x"3400";
            when "11" & x"947" => DATA <= x"10a0";
            when "11" & x"948" => DATA <= x"0080";
            when "11" & x"949" => DATA <= x"0041";
            when "11" & x"94a" => DATA <= x"400a";
            when "11" & x"94b" => DATA <= x"2010";
            when "11" & x"94c" => DATA <= x"8bc0";
            when "11" & x"94d" => DATA <= x"3400";
            when "11" & x"94e" => DATA <= x"4000";
            when "11" & x"94f" => DATA <= x"1000";
            when "11" & x"950" => DATA <= x"041e";
            when "11" & x"951" => DATA <= x"0020";
            when "11" & x"952" => DATA <= x"f00f";
            when "11" & x"953" => DATA <= x"0000";
            when "11" & x"954" => DATA <= x"00bc";
            when "11" & x"955" => DATA <= x"02c0";
            when "11" & x"956" => DATA <= x"0434";
            when "11" & x"957" => DATA <= x"0003";
            when "11" & x"958" => DATA <= x"a001";
            when "11" & x"959" => DATA <= x"4a02";
            when "11" & x"95a" => DATA <= x"8001";
            when "11" & x"95b" => DATA <= x"1e00";
            when "11" & x"95c" => DATA <= x"0020";
            when "11" & x"95d" => DATA <= x"7800";
            when "11" & x"95e" => DATA <= x"0821";
            when "11" & x"95f" => DATA <= x"4007";
            when "11" & x"960" => DATA <= x"aa00";
            when "11" & x"961" => DATA <= x"0848";
            when "11" & x"962" => DATA <= x"03ff";
            when "11" & x"963" => DATA <= x"c01f";
            when "11" & x"964" => DATA <= x"fe00";
            when "11" & x"965" => DATA <= x"fff0";
            when "11" & x"966" => DATA <= x"01fd";
            when "11" & x"967" => DATA <= x"0004";
            when "11" & x"968" => DATA <= x"3c03";
            when "11" & x"969" => DATA <= x"4004";
            when "11" & x"96a" => DATA <= x"1200";
            when "11" & x"96b" => DATA <= x"10a0";
            when "11" & x"96c" => DATA <= x"0085";
            when "11" & x"96d" => DATA <= x"0004";
            when "11" & x"96e" => DATA <= x"3c03";
            when "11" & x"96f" => DATA <= x"4010";
            when "11" & x"970" => DATA <= x"1e00";
            when "11" & x"971" => DATA <= x"fff0";
            when "11" & x"972" => DATA <= x"07bf";
            when "11" & x"973" => DATA <= x"803e";
            when "11" & x"974" => DATA <= x"ec00";
            when "11" & x"975" => DATA <= x"c005";
            when "11" & x"976" => DATA <= x"a001";
            when "11" & x"977" => DATA <= x"0700";
            when "11" & x"978" => DATA <= x"007c";
            when "11" & x"979" => DATA <= x"02c0";
            when "11" & x"97a" => DATA <= x"0600";
            when "11" & x"97b" => DATA <= x"0300";
            when "11" & x"97c" => DATA <= x"0041";
            when "11" & x"97d" => DATA <= x"e014";
            when "11" & x"97e" => DATA <= x"0040";
            when "11" & x"97f" => DATA <= x"9000";
            when "11" & x"980" => DATA <= x"8700";
            when "11" & x"981" => DATA <= x"0801";
            when "11" & x"982" => DATA <= x"1400";
            when "11" & x"983" => DATA <= x"08e0";
            when "11" & x"984" => DATA <= x"006d";
            when "11" & x"985" => DATA <= x"0020";
            when "11" & x"986" => DATA <= x"3c03";
            when "11" & x"987" => DATA <= x"c03c";
            when "11" & x"988" => DATA <= x"0280";
            when "11" & x"989" => DATA <= x"041e";
            when "11" & x"98a" => DATA <= x"0020";
            when "11" & x"98b" => DATA <= x"0c70";
            when "11" & x"98c" => DATA <= x"0004";
            when "11" & x"98d" => DATA <= x"4160";
            when "11" & x"98e" => DATA <= x"0200";
            when "11" & x"98f" => DATA <= x"0800";
            when "11" & x"990" => DATA <= x"1140";
            when "11" & x"991" => DATA <= x"0080";
            when "11" & x"992" => DATA <= x"0004";
            when "11" & x"993" => DATA <= x"3c00";
            when "11" & x"994" => DATA <= x"a0ef";
            when "11" & x"995" => DATA <= x"00d0";
            when "11" & x"996" => DATA <= x"0040";
            when "11" & x"997" => DATA <= x"0141";
            when "11" & x"998" => DATA <= x"a00e";
            when "11" & x"999" => DATA <= x"c7e3";
            when "11" & x"99a" => DATA <= x"e1d8";
            when "11" & x"99b" => DATA <= x"fc7c";
            when "11" & x"99c" => DATA <= x"3f9f";
            when "11" & x"99d" => DATA <= x"167e";
            when "11" & x"99e" => DATA <= x"bf1f";
            when "11" & x"99f" => DATA <= x"d7f8";
            when "11" & x"9a0" => DATA <= x"02bf";
            when "11" & x"9a1" => DATA <= x"8015";
            when "11" & x"9a2" => DATA <= x"fe2b";
            when "11" & x"9a3" => DATA <= x"1780";
            when "11" & x"9a4" => DATA <= x"0560";
            when "11" & x"9a5" => DATA <= x"a200";
            when "11" & x"9a6" => DATA <= x"b42e";
            when "11" & x"9a7" => DATA <= x"01b0";
            when "11" & x"9a8" => DATA <= x"0482";
            when "11" & x"9a9" => DATA <= x"2900";
            when "11" & x"9aa" => DATA <= x"8b44";
            when "11" & x"9ab" => DATA <= x"a210";
            when "11" & x"9ac" => DATA <= x"08a5";
            when "11" & x"9ad" => DATA <= x"51fc";
            when "11" & x"9ae" => DATA <= x"8f4f";
            when "11" & x"9af" => DATA <= x"effa";
            when "11" & x"9b0" => DATA <= x"7f23";
            when "11" & x"9b1" => DATA <= x"be00";
            when "11" & x"9b2" => DATA <= x"5400";
            when "11" & x"9b3" => DATA <= x"fb00";
            when "11" & x"9b4" => DATA <= x"0200";
            when "11" & x"9b5" => DATA <= x"4ffe";
            when "11" & x"9b6" => DATA <= x"0001";
            when "11" & x"9b7" => DATA <= x"f000";
            when "11" & x"9b8" => DATA <= x"fdc0";
            when "11" & x"9b9" => DATA <= x"0098";
            when "11" & x"9ba" => DATA <= x"0702";
            when "11" & x"9bb" => DATA <= x"001f";
            when "11" & x"9bc" => DATA <= x"7ffd";
            when "11" & x"9bd" => DATA <= x"e6fb";
            when "11" & x"9be" => DATA <= x"eff7";
            when "11" & x"9bf" => DATA <= x"df80";
            when "11" & x"9c0" => DATA <= x"847c";
            when "11" & x"9c1" => DATA <= x"0000";
            when "11" & x"9c2" => DATA <= x"e777";
            when "11" & x"9c3" => DATA <= x"b9e7";
            when "11" & x"9c4" => DATA <= x"bdfe";
            when "11" & x"9c5" => DATA <= x"805c";
            when "11" & x"9c6" => DATA <= x"0eb6";
            when "11" & x"9c7" => DATA <= x"fb40";
            when "11" & x"9c8" => DATA <= x"2bfc";
            when "11" & x"9c9" => DATA <= x"1fa0";
            when "11" & x"9ca" => DATA <= x"0ff6";
            when "11" & x"9cb" => DATA <= x"0380";
            when "11" & x"9cc" => DATA <= x"00e0";
            when "11" & x"9cd" => DATA <= x"7130";
            when "11" & x"9ce" => DATA <= x"9c0c";
            when "11" & x"9cf" => DATA <= x"0703";
            when "11" & x"9d0" => DATA <= x"8e87";
            when "11" & x"9d1" => DATA <= x"d3f4";
            when "11" & x"9d2" => DATA <= x"3e1e";
            when "11" & x"9d3" => DATA <= x"09a7";
            when "11" & x"9d4" => DATA <= x"c2b4";
            when "11" & x"9d5" => DATA <= x"0a0d";
            when "11" & x"9d6" => DATA <= x"0050";
            when "11" & x"9d7" => DATA <= x"2014";
            when "11" & x"9d8" => DATA <= x"fc54";
            when "11" & x"9d9" => DATA <= x"0017";
            when "11" & x"9da" => DATA <= x"c21c";
            when "11" & x"9db" => DATA <= x"a9bf";
            when "11" & x"9dc" => DATA <= x"d5fe";
            when "11" & x"9dd" => DATA <= x"fe00";
            when "11" & x"9de" => DATA <= x"d000";
            when "11" & x"9df" => DATA <= x"4000";
            when "11" & x"9e0" => DATA <= x"b8d0";
            when "11" & x"9e1" => DATA <= x"0040";
            when "11" & x"9e2" => DATA <= x"01bf";
            when "11" & x"9e3" => DATA <= x"e00e";
            when "11" & x"9e4" => DATA <= x"fa00";
            when "11" & x"9e5" => DATA <= x"1048";
            when "11" & x"9e6" => DATA <= x"01fa";
            when "11" & x"9e7" => DATA <= x"8002";
            when "11" & x"9e8" => DATA <= x"1400";
            when "11" & x"9e9" => DATA <= x"0200";
            when "11" & x"9ea" => DATA <= x"2df4";
            when "11" & x"9eb" => DATA <= x"0102";
            when "11" & x"9ec" => DATA <= x"006d";
            when "11" & x"9ed" => DATA <= x"e801";
            when "11" & x"9ee" => DATA <= x"0000";
            when "11" & x"9ef" => DATA <= x"edf0";
            when "11" & x"9f0" => DATA <= x"03f7";
            when "11" & x"9f1" => DATA <= x"8006";
            when "11" & x"9f2" => DATA <= x"fc03";
            when "11" & x"9f3" => DATA <= x"c024";
            when "11" & x"9f4" => DATA <= x"0021";
            when "11" & x"9f5" => DATA <= x"a001";
            when "11" & x"9f6" => DATA <= x"0031";
            when "11" & x"9f7" => DATA <= x"0280";
            when "11" & x"9f8" => DATA <= x"009c";
            when "11" & x"9f9" => DATA <= x"0080";
            when "11" & x"9fa" => DATA <= x"0878";
            when "11" & x"9fb" => DATA <= x"0780";
            when "11" & x"9fc" => DATA <= x"5800";
            when "11" & x"9fd" => DATA <= x"4280";
            when "11" & x"9fe" => DATA <= x"0412";
            when "11" & x"9ff" => DATA <= x"0020";
            when "11" & x"a00" => DATA <= x"0008";
            when "11" & x"a01" => DATA <= x"b801";
            when "11" & x"a02" => DATA <= x"01c0";
            when "11" & x"a03" => DATA <= x"001f";
            when "11" & x"a04" => DATA <= x"00f0";
            when "11" & x"a05" => DATA <= x"0000";
            when "11" & x"a06" => DATA <= x"07c0";
            when "11" & x"a07" => DATA <= x"3803";
            when "11" & x"a08" => DATA <= x"80bc";
            when "11" & x"a09" => DATA <= x"02c0";
            when "11" & x"a0a" => DATA <= x"1012";
            when "11" & x"a0b" => DATA <= x"0008";
            when "11" & x"a0c" => DATA <= x"1500";
            when "11" & x"a0d" => DATA <= x"1008";
            when "11" & x"a0e" => DATA <= x"221a";
            when "11" & x"a0f" => DATA <= x"0000";
            when "11" & x"a10" => DATA <= x"61f0";
            when "11" & x"a11" => DATA <= x"0e00";
            when "11" & x"a12" => DATA <= x"0168";
            when "11" & x"a13" => DATA <= x"000a";
            when "11" & x"a14" => DATA <= x"8004";
            when "11" & x"a15" => DATA <= x"6001";
            when "11" & x"a16" => DATA <= x"d800";
            when "11" & x"a17" => DATA <= x"05c0";
            when "11" & x"a18" => DATA <= x"0100";
            when "11" & x"a19" => DATA <= x"0282";
            when "11" & x"a1a" => DATA <= x"8010";
            when "11" & x"a1b" => DATA <= x"3400";
            when "11" & x"a1c" => DATA <= x"0800";
            when "11" & x"a1d" => DATA <= x"0228";
            when "11" & x"a1e" => DATA <= x"0081";
            when "11" & x"a1f" => DATA <= x"2008";
            when "11" & x"a20" => DATA <= x"da00";
            when "11" & x"a21" => DATA <= x"1050";
            when "11" & x"a22" => DATA <= x"0010";
            when "11" & x"a23" => DATA <= x"000c";
            when "11" & x"a24" => DATA <= x"f00f";
            when "11" & x"a25" => DATA <= x"00b0";
            when "11" & x"a26" => DATA <= x"0085";
            when "11" & x"a27" => DATA <= x"0004";
            when "11" & x"a28" => DATA <= x"2400";
            when "11" & x"a29" => DATA <= x"41c0";
            when "11" & x"a2a" => DATA <= x"010b";
            when "11" & x"a2b" => DATA <= x"0040";
            when "11" & x"a2c" => DATA <= x"6800";
            when "11" & x"a2d" => DATA <= x"1000";
            when "11" & x"a2e" => DATA <= x"66d0";
            when "11" & x"a2f" => DATA <= x"0010";
            when "11" & x"a30" => DATA <= x"0029";
            when "11" & x"a31" => DATA <= x"4001";
            when "11" & x"a32" => DATA <= x"0a00";
            when "11" & x"a33" => DATA <= x"4080";
            when "11" & x"a34" => DATA <= x"1154";
            when "11" & x"a35" => DATA <= x"0018";
            when "11" & x"a36" => DATA <= x"0810";
            when "11" & x"a37" => DATA <= x"0e00";
            when "11" & x"a38" => DATA <= x"0381";
            when "11" & x"a39" => DATA <= x"40e1";
            when "11" & x"a3a" => DATA <= x"c000";
            when "11" & x"a3b" => DATA <= x"1000";
            when "11" & x"a3c" => DATA <= x"0400";
            when "11" & x"a3d" => DATA <= x"01e0";
            when "11" & x"a3e" => DATA <= x"0027";
            when "11" & x"a3f" => DATA <= x"8050";
            when "11" & x"a40" => DATA <= x"000c";
            when "11" & x"a41" => DATA <= x"0200";
            when "11" & x"a42" => DATA <= x"2150";
            when "11" & x"a43" => DATA <= x"0108";
            when "11" & x"a44" => DATA <= x"01c0";
            when "11" & x"a45" => DATA <= x"440e";
            when "11" & x"a46" => DATA <= x"0008";
            when "11" & x"a47" => DATA <= x"6800";
            when "11" & x"a48" => DATA <= x"2340";
            when "11" & x"a49" => DATA <= x"0080";
            when "11" & x"a4a" => DATA <= x"0085";
            when "11" & x"a4b" => DATA <= x"4050";
            when "11" & x"a4c" => DATA <= x"0202";
            when "11" & x"a4d" => DATA <= x"4008";
            when "11" & x"a4e" => DATA <= x"1400";
            when "11" & x"a4f" => DATA <= x"f0a0";
            when "11" & x"a50" => DATA <= x"0024";
            when "11" & x"a51" => DATA <= x"8030";
            when "11" & x"a52" => DATA <= x"0056";
            when "11" & x"a53" => DATA <= x"0029";
            when "11" & x"a54" => DATA <= x"d000";
            when "11" & x"a55" => DATA <= x"8000";
            when "11" & x"a56" => DATA <= x"4140";
            when "11" & x"a57" => DATA <= x"021f";
            when "11" & x"a58" => DATA <= x"0000";
            when "11" & x"a59" => DATA <= x"8001";
            when "11" & x"a5a" => DATA <= x"0010";
            when "11" & x"a5b" => DATA <= x"0063";
            when "11" & x"a5c" => DATA <= x"c008";
            when "11" & x"a5d" => DATA <= x"1e00";
            when "11" & x"a5e" => DATA <= x"0014";
            when "11" & x"a5f" => DATA <= x"2201";
            when "11" & x"a60" => DATA <= x"0007";
            when "11" & x"a61" => DATA <= x"c700";
            when "11" & x"a62" => DATA <= x"3e1f";
            when "11" & x"a63" => DATA <= x"ce87";
            when "11" & x"a64" => DATA <= x"c3fd";
            when "11" & x"a65" => DATA <= x"d8fc";
            when "11" & x"a66" => DATA <= x"7c51";
            when "11" & x"a67" => DATA <= x"fd5f";
            when "11" & x"a68" => DATA <= x"d1fa";
            when "11" & x"a69" => DATA <= x"fc7f";
            when "11" & x"a6a" => DATA <= x"4015";
            when "11" & x"a6b" => DATA <= x"fe00";
            when "11" & x"a6c" => DATA <= x"7f9f";
            when "11" & x"a6d" => DATA <= x"c001";
            when "11" & x"a6e" => DATA <= x"c005";
            when "11" & x"a6f" => DATA <= x"0300";
            when "11" & x"a70" => DATA <= x"0034";
            when "11" & x"a71" => DATA <= x"015e";
            when "11" & x"a72" => DATA <= x"0e0a";
            when "11" & x"a73" => DATA <= x"f048";
            when "11" & x"a74" => DATA <= x"001e";
            when "11" & x"a75" => DATA <= x"0a8a";
            when "11" & x"a76" => DATA <= x"aa51";
            when "11" & x"a77" => DATA <= x"2090";
            when "11" & x"a78" => DATA <= x"08a7";
            when "11" & x"a79" => DATA <= x"57bf";
            when "11" & x"a7a" => DATA <= x"9fdf";
            when "11" & x"a7b" => DATA <= x"8b80";
            when "11" & x"a7c" => DATA <= x"c305";
            when "11" & x"a7d" => DATA <= x"8b40";
            when "11" & x"a7e" => DATA <= x"0227";
            when "11" & x"a7f" => DATA <= x"fb84";
            when "11" & x"a80" => DATA <= x"0007";
            when "11" & x"a81" => DATA <= x"7fbf";
            when "11" & x"a82" => DATA <= x"0000";
            when "11" & x"a83" => DATA <= x"4aff";
            when "11" & x"a84" => DATA <= x"7800";
            when "11" & x"a85" => DATA <= x"01e0";
            when "11" & x"a86" => DATA <= x"1a80";
            when "11" & x"a87" => DATA <= x"eff6";
            when "11" & x"a88" => DATA <= x"0001";
            when "11" & x"a89" => DATA <= x"800f";
            when "11" & x"a8a" => DATA <= x"3ff7";
            when "11" & x"a8b" => DATA <= x"fbed";
            when "11" & x"a8c" => DATA <= x"e0e3";
            when "11" & x"a8d" => DATA <= x"5934";
            when "11" & x"a8e" => DATA <= x"e5c6";
            when "11" & x"a8f" => DATA <= x"4040";
            when "11" & x"a90" => DATA <= x"010b";
            when "11" & x"a91" => DATA <= x"007f";
            when "11" & x"a92" => DATA <= x"bbcd";
            when "11" & x"a93" => DATA <= x"e077";
            when "11" & x"a94" => DATA <= x"3abd";
            when "11" & x"a95" => DATA <= x"daef";
            when "11" & x"a96" => DATA <= x"1f80";
            when "11" & x"a97" => DATA <= x"8000";
            when "11" & x"a98" => DATA <= x"2000";
            when "11" & x"a99" => DATA <= x"a86c";
            when "11" & x"a9a" => DATA <= x"3e00";
            when "11" & x"a9b" => DATA <= x"3c2c";
            when "11" & x"a9c" => DATA <= x"01f8";
            when "11" & x"a9d" => DATA <= x"ffb0";
            when "11" & x"a9e" => DATA <= x"073b";
            when "11" & x"a9f" => DATA <= x"3dcc";
            when "11" & x"aa0" => DATA <= x"02ae";
            when "11" & x"aa1" => DATA <= x"0603";
            when "11" & x"aa2" => DATA <= x"f836";
            when "11" & x"aa3" => DATA <= x"1f4f";
            when "11" & x"aa4" => DATA <= x"83c3";
            when "11" & x"aa5" => DATA <= x"e9f0";
            when "11" & x"aa6" => DATA <= x"fa7c";
            when "11" & x"aa7" => DATA <= x"0800";
            when "11" & x"aa8" => DATA <= x"0201";
            when "11" & x"aa9" => DATA <= x"7804";
            when "11" & x"aaa" => DATA <= x"0800";
            when "11" & x"aab" => DATA <= x"2a10";
            when "11" & x"aac" => DATA <= x"0000";
            when "11" & x"aad" => DATA <= x"40a0";
            when "11" & x"aae" => DATA <= x"00ab";
            when "11" & x"aaf" => DATA <= x"dfc7";
            when "11" & x"ab0" => DATA <= x"eefe";
            when "11" & x"ab1" => DATA <= x"7fbe";
            when "11" & x"ab2" => DATA <= x"2400";
            when "11" & x"ab3" => DATA <= x"0200";
            when "11" & x"ab4" => DATA <= x"5c37";
            when "11" & x"ab5" => DATA <= x"6c01";
            when "11" & x"ab6" => DATA <= x"aabf";
            when "11" & x"ab7" => DATA <= x"e000";
            when "11" & x"ab8" => DATA <= x"1500";
            when "11" & x"ab9" => DATA <= x"3fcd";
            when "11" & x"aba" => DATA <= x"b600";
            when "11" & x"abb" => DATA <= x"ef5f";
            when "11" & x"abc" => DATA <= x"f000";
            when "11" & x"abd" => DATA <= x"1280";
            when "11" & x"abe" => DATA <= x"16ef";
            when "11" & x"abf" => DATA <= x"bb00";
            when "11" & x"ac0" => DATA <= x"6dbf";
            when "11" & x"ac1" => DATA <= x"6c01";
            when "11" & x"ac2" => DATA <= x"fa4e";
            when "11" & x"ac3" => DATA <= x"b007";
            when "11" & x"ac4" => DATA <= x"f846";
            when "11" & x"ac5" => DATA <= x"8002";
            when "11" & x"ac6" => DATA <= x"014a";
            when "11" & x"ac7" => DATA <= x"001f";
            when "11" & x"ac8" => DATA <= x"f000";
            when "11" & x"ac9" => DATA <= x"07c0";
            when "11" & x"aca" => DATA <= x"041a";
            when "11" & x"acb" => DATA <= x"0010";
            when "11" & x"acc" => DATA <= x"0308";
            when "11" & x"acd" => DATA <= x"3800";
            when "11" & x"ace" => DATA <= x"09a0";
            when "11" & x"acf" => DATA <= x"040f";
            when "11" & x"ad0" => DATA <= x"00f0";
            when "11" & x"ad1" => DATA <= x"0900";
            when "11" & x"ad2" => DATA <= x"0850";
            when "11" & x"ad3" => DATA <= x"0043";
            when "11" & x"ad4" => DATA <= x"8002";
            when "11" & x"ad5" => DATA <= x"2200";
            when "11" & x"ad6" => DATA <= x"008a";
            when "11" & x"ad7" => DATA <= x"8004";
            when "11" & x"ad8" => DATA <= x"1e01";
            when "11" & x"ad9" => DATA <= x"6003";
            when "11" & x"ada" => DATA <= x"0f00";
            when "11" & x"adb" => DATA <= x"f00b";
            when "11" & x"adc" => DATA <= x"0001";
            when "11" & x"add" => DATA <= x"5000";
            when "11" & x"ade" => DATA <= x"4804";
            when "11" & x"adf" => DATA <= x"00a0";
            when "11" & x"ae0" => DATA <= x"2f00";
            when "11" & x"ae1" => DATA <= x"a001";
            when "11" & x"ae2" => DATA <= x"0d80";
            when "11" & x"ae3" => DATA <= x"2000";
            when "11" & x"ae4" => DATA <= x"1500";
            when "11" & x"ae5" => DATA <= x"0060";
            when "11" & x"ae6" => DATA <= x"1011";
            when "11" & x"ae7" => DATA <= x"0002";
            when "11" & x"ae8" => DATA <= x"0580";
            when "11" & x"ae9" => DATA <= x"2000";
            when "11" & x"aea" => DATA <= x"1501";
            when "11" & x"aeb" => DATA <= x"c00c";
            when "11" & x"aec" => DATA <= x"27dd";
            when "11" & x"aed" => DATA <= x"0004";
            when "11" & x"aee" => DATA <= x"4000";
            when "11" & x"aef" => DATA <= x"2000";
            when "11" & x"af0" => DATA <= x"45ff";
            when "11" & x"af1" => DATA <= x"e00f";
            when "11" & x"af2" => DATA <= x"ef00";
            when "11" & x"af3" => DATA <= x"7ff8";
            when "11" & x"af4" => DATA <= x"00ff";
            when "11" & x"af5" => DATA <= x"c03c";
            when "11" & x"af6" => DATA <= x"0000";
            when "11" & x"af7" => DATA <= x"20f0";
            when "11" & x"af8" => DATA <= x"0085";
            when "11" & x"af9" => DATA <= x"0004";
            when "11" & x"afa" => DATA <= x"3802";
            when "11" & x"afb" => DATA <= x"8428";
            when "11" & x"afc" => DATA <= x"0021";
            when "11" & x"afd" => DATA <= x"c001";
            when "11" & x"afe" => DATA <= x"1407";
            when "11" & x"aff" => DATA <= x"803b";
            when "11" & x"b00" => DATA <= x"fc01";
            when "11" & x"b01" => DATA <= x"efe0";
            when "11" & x"b02" => DATA <= x"0fff";
            when "11" & x"b03" => DATA <= x"003b";
            when "11" & x"b04" => DATA <= x"8001";
            when "11" & x"b05" => DATA <= x"0100";
            when "11" & x"b06" => DATA <= x"0102";
            when "11" & x"b07" => DATA <= x"8000";
            when "11" & x"b08" => DATA <= x"3e01";
            when "11" & x"b09" => DATA <= x"e000";
            when "11" & x"b0a" => DATA <= x"0012";
            when "11" & x"b0b" => DATA <= x"0000";
            when "11" & x"b0c" => DATA <= x"0640";
            when "11" & x"b0d" => DATA <= x"5000";
            when "11" & x"b0e" => DATA <= x"0404";
            when "11" & x"b0f" => DATA <= x"0001";
            when "11" & x"b10" => DATA <= x"1080";
            when "11" & x"b11" => DATA <= x"0420";
            when "11" & x"b12" => DATA <= x"0008";
            when "11" & x"b13" => DATA <= x"21a0";
            when "11" & x"b14" => DATA <= x"010f";
            when "11" & x"b15" => DATA <= x"0000";
            when "11" & x"b16" => DATA <= x"0228";
            when "11" & x"b17" => DATA <= x"0009";
            when "11" & x"b18" => DATA <= x"4000";
            when "11" & x"b19" => DATA <= x"4200";
            when "11" & x"b1a" => DATA <= x"6240";
            when "11" & x"b1b" => DATA <= x"1c06";
            when "11" & x"b1c" => DATA <= x"0183";
            when "11" & x"b1d" => DATA <= x"c240";
            when "11" & x"b1e" => DATA <= x"0805";
            when "11" & x"b1f" => DATA <= x"e401";
            when "11" & x"b20" => DATA <= x"4340";
            when "11" & x"b21" => DATA <= x"0060";
            when "11" & x"b22" => DATA <= x"1000";
            when "11" & x"b23" => DATA <= x"6380";
            when "11" & x"b24" => DATA <= x"003e";
            when "11" & x"b25" => DATA <= x"0001";
            when "11" & x"b26" => DATA <= x"a001";
            when "11" & x"b27" => DATA <= x"0c80";
            when "11" & x"b28" => DATA <= x"0068";
            when "11" & x"b29" => DATA <= x"0002";
            when "11" & x"b2a" => DATA <= x"6190";
            when "11" & x"b2b" => DATA <= x"0100";
            when "11" & x"b2c" => DATA <= x"00c9";
            when "11" & x"b2d" => DATA <= x"a000";
            when "11" & x"b2e" => DATA <= x"8b00";
            when "11" & x"b2f" => DATA <= x"a085";
            when "11" & x"b30" => DATA <= x"4021";
            when "11" & x"b31" => DATA <= x"fcfc";
            when "11" & x"b32" => DATA <= x"7c3f";
            when "11" & x"b33" => DATA <= x"abe1";
            when "11" & x"b34" => DATA <= x"fce8";
            when "11" & x"b35" => DATA <= x"e3f5";
            when "11" & x"b36" => DATA <= x"ff1f";
            when "11" & x"b37" => DATA <= x"afd7";
            when "11" & x"b38" => DATA <= x"cbf0";
            when "11" & x"b39" => DATA <= x"027c";
            when "11" & x"b3a" => DATA <= x"bf48";
            when "11" & x"b3b" => DATA <= x"03f0";
            when "11" & x"b3c" => DATA <= x"2228";
            when "11" & x"b3d" => DATA <= x"6140";
            when "11" & x"b3e" => DATA <= x"0161";
            when "11" & x"b3f" => DATA <= x"0098";
            when "11" & x"b40" => DATA <= x"0010";
            when "11" & x"b41" => DATA <= x"6380";
            when "11" & x"b42" => DATA <= x"1800";
            when "11" & x"b43" => DATA <= x"0600";
            when "11" & x"b44" => DATA <= x"0110";
            when "11" & x"b45" => DATA <= x"8a61";
            when "11" & x"b46" => DATA <= x"2290";
            when "11" & x"b47" => DATA <= x"2825";
            when "11" & x"b48" => DATA <= x"42aa";
            when "11" & x"b49" => DATA <= x"5fcd";
            when "11" & x"b4a" => DATA <= x"fcfe";
            when "11" & x"b4b" => DATA <= x"0002";
            when "11" & x"b4c" => DATA <= x"7003";
            when "11" & x"b4d" => DATA <= x"1402";
            when "11" & x"b4e" => DATA <= x"f8a0";
            when "11" & x"b4f" => DATA <= x"0020";
            when "11" & x"b50" => DATA <= x"01f8";
            when "11" & x"b51" => DATA <= x"ff90";
            when "11" & x"b52" => DATA <= x"0a80";
            when "11" & x"b53" => DATA <= x"40d4";
            when "11" & x"b54" => DATA <= x"7b83";
            when "11" & x"b55" => DATA <= x"ffeb";
            when "11" & x"b56" => DATA <= x"febe";
            when "11" & x"b57" => DATA <= x"dfef";
            when "11" & x"b58" => DATA <= x"beff";
            when "11" & x"b59" => DATA <= x"0048";
            when "11" & x"b5a" => DATA <= x"0f38";
            when "11" & x"b5b" => DATA <= x"e800";
            when "11" & x"b5c" => DATA <= x"4280";
            when "11" & x"b5d" => DATA <= x"1df3";
            when "11" & x"b5e" => DATA <= x"feef";
            when "11" & x"b5f" => DATA <= x"03b9";
            when "11" & x"b60" => DATA <= x"e8f9";
            when "11" & x"b61" => DATA <= x"7cbf";
            when "11" & x"b62" => DATA <= x"07d0";
            when "11" & x"b63" => DATA <= x"0081";
            when "11" & x"b64" => DATA <= x"f87c";
            when "11" & x"b65" => DATA <= x"2780";
            when "11" & x"b66" => DATA <= x"5c1c";
            when "11" & x"b67" => DATA <= x"00ff";
            when "11" & x"b68" => DATA <= x"603c";
            when "11" & x"b69" => DATA <= x"0f8f";
            when "11" & x"b6a" => DATA <= x"fe00";
            when "11" & x"b6b" => DATA <= x"77b0";
            when "11" & x"b6c" => DATA <= x"dcfd";
            when "11" & x"b6d" => DATA <= x"c000";
            when "11" & x"b6e" => DATA <= x"7107";
            when "11" & x"b6f" => DATA <= x"c369";
            when "11" & x"b70" => DATA <= x"f0f8";
            when "11" & x"b71" => DATA <= x"7b87";
            when "11" & x"b72" => DATA <= x"c000";
            when "11" & x"b73" => DATA <= x"412d";
            when "11" & x"b74" => DATA <= x"0200";
            when "11" & x"b75" => DATA <= x"2914";
            when "11" & x"b76" => DATA <= x"2940";
            when "11" & x"b77" => DATA <= x"054a";
            when "11" & x"b78" => DATA <= x"002a";
            when "11" & x"b79" => DATA <= x"143b";
            when "11" & x"b7a" => DATA <= x"f9ff";
            when "11" & x"b7b" => DATA <= x"3fc1";
            when "11" & x"b7c" => DATA <= x"0002";
            when "11" & x"b7d" => DATA <= x"e280";
            when "11" & x"b7e" => DATA <= x"1514";
            when "11" & x"b7f" => DATA <= x"0008";
            when "11" & x"b80" => DATA <= x"0037";
            when "11" & x"b81" => DATA <= x"e800";
            when "11" & x"b82" => DATA <= x"8400";
            when "11" & x"b83" => DATA <= x"40d0";
            when "11" & x"b84" => DATA <= x"03fe";
            when "11" & x"b85" => DATA <= x"8017";
            when "11" & x"b86" => DATA <= x"6002";
            when "11" & x"b87" => DATA <= x"0500";
            when "11" & x"b88" => DATA <= x"1fe8";
            when "11" & x"b89" => DATA <= x"00a0";
            when "11" & x"b8a" => DATA <= x"0010";
            when "11" & x"b8b" => DATA <= x"5002";
            when "11" & x"b8c" => DATA <= x"fe80";
            when "11" & x"b8d" => DATA <= x"0114";
            when "11" & x"b8e" => DATA <= x"0081";
            when "11" & x"b8f" => DATA <= x"0036";
            when "11" & x"b90" => DATA <= x"f400";
            when "11" & x"b91" => DATA <= x"8000";
            when "11" & x"b92" => DATA <= x"7ed0";
            when "11" & x"b93" => DATA <= x"0282";
            when "11" & x"b94" => DATA <= x"400d";
            when "11" & x"b95" => DATA <= x"d400";
            when "11" & x"b96" => DATA <= x"4a00";
            when "11" & x"b97" => DATA <= x"0128";
            when "11" & x"b98" => DATA <= x"0037";
            when "11" & x"b99" => DATA <= x"4001";
            when "11" & x"b9a" => DATA <= x"1000";
            when "11" & x"b9b" => DATA <= x"0bc0";
            when "11" & x"b9c" => DATA <= x"3c02";
            when "11" & x"b9d" => DATA <= x"8000";
            when "11" & x"b9e" => DATA <= x"400a";
            when "11" & x"b9f" => DATA <= x"011b";
            when "11" & x"ba0" => DATA <= x"8000";
            when "11" & x"ba1" => DATA <= x"21fe";
            when "11" & x"ba2" => DATA <= x"0001";
            when "11" & x"ba3" => DATA <= x"7002";
            when "11" & x"ba4" => DATA <= x"03c0";
            when "11" & x"ba5" => DATA <= x"021e";
            when "11" & x"ba6" => DATA <= x"01c0";
            when "11" & x"ba7" => DATA <= x"010a";
            when "11" & x"ba8" => DATA <= x"0008";
            when "11" & x"ba9" => DATA <= x"4800";
            when "11" & x"baa" => DATA <= x"8804";
            when "11" & x"bab" => DATA <= x"2210";
            when "11" & x"bac" => DATA <= x"0084";
            when "11" & x"bad" => DATA <= x"480f";
            when "11" & x"bae" => DATA <= x"00e0";
            when "11" & x"baf" => DATA <= x"0107";
            when "11" & x"bb0" => DATA <= x"0020";
            when "11" & x"bb1" => DATA <= x"2400";
            when "11" & x"bb2" => DATA <= x"0340";
            when "11" & x"bb3" => DATA <= x"001f";
            when "11" & x"bb4" => DATA <= x"0000";
            when "11" & x"bb5" => DATA <= x"0080";
            when "11" & x"bb6" => DATA <= x"002f";
            when "11" & x"bb7" => DATA <= x"0000";
            when "11" & x"bb8" => DATA <= x"0078";
            when "11" & x"bb9" => DATA <= x"0011";
            when "11" & x"bba" => DATA <= x"c002";
            when "11" & x"bbb" => DATA <= x"0040";
            when "11" & x"bbc" => DATA <= x"0042";
            when "11" & x"bbd" => DATA <= x"0060";
            when "11" & x"bbe" => DATA <= x"101c";
            when "11" & x"bbf" => DATA <= x"0003";
            when "11" & x"bc0" => DATA <= x"4d00";
            when "11" & x"bc1" => DATA <= x"30ec";
            when "11" & x"bc2" => DATA <= x"0080";
            when "11" & x"bc3" => DATA <= x"0060";
            when "11" & x"bc4" => DATA <= x"001c";
            when "11" & x"bc5" => DATA <= x"1200";
            when "11" & x"bc6" => DATA <= x"f001";
            when "11" & x"bc7" => DATA <= x"800f";
            when "11" & x"bc8" => DATA <= x"7400";
            when "11" & x"bc9" => DATA <= x"f000";
            when "11" & x"bca" => DATA <= x"00e8";
            when "11" & x"bcb" => DATA <= x"0163";
            when "11" & x"bcc" => DATA <= x"400b";
            when "11" & x"bcd" => DATA <= x"7a00";
            when "11" & x"bce" => DATA <= x"0400";
            when "11" & x"bcf" => DATA <= x"1b34";
            when "11" & x"bd0" => DATA <= x"0057";
            when "11" & x"bd1" => DATA <= x"0020";
            when "11" & x"bd2" => DATA <= x"6801";
            when "11" & x"bd3" => DATA <= x"db40";
            when "11" & x"bd4" => DATA <= x"0bd0";
            when "11" & x"bd5" => DATA <= x"0100";
            when "11" & x"bd6" => DATA <= x"0800";
            when "11" & x"bd7" => DATA <= x"1750";
            when "11" & x"bd8" => DATA <= x"006c";
            when "11" & x"bd9" => DATA <= x"0020";
            when "11" & x"bda" => DATA <= x"f00e";
            when "11" & x"bdb" => DATA <= x"0010";
            when "11" & x"bdc" => DATA <= x"7800";
            when "11" & x"bdd" => DATA <= x"43c0";
            when "11" & x"bde" => DATA <= x"2442";
            when "11" & x"bdf" => DATA <= x"4010";
            when "11" & x"be0" => DATA <= x"1400";
            when "11" & x"be1" => DATA <= x"8000";
            when "11" & x"be2" => DATA <= x"1000";
            when "11" & x"be3" => DATA <= x"8003";
            when "11" & x"be4" => DATA <= x"7500";
            when "11" & x"be5" => DATA <= x"3bc0";
            when "11" & x"be6" => DATA <= x"0200";
            when "11" & x"be7" => DATA <= x"1001";
            when "11" & x"be8" => DATA <= x"6f40";
            when "11" & x"be9" => DATA <= x"0ff0";
            when "11" & x"bea" => DATA <= x"0080";
            when "11" & x"beb" => DATA <= x"0200";
            when "11" & x"bec" => DATA <= x"4dd0";
            when "11" & x"bed" => DATA <= x"03b8";
            when "11" & x"bee" => DATA <= x"0010";
            when "11" & x"bef" => DATA <= x"3800";
            when "11" & x"bf0" => DATA <= x"0f25";
            when "11" & x"bf1" => DATA <= x"0381";
            when "11" & x"bf2" => DATA <= x"5400";
            when "11" & x"bf3" => DATA <= x"7800";
            when "11" & x"bf4" => DATA <= x"8000";
            when "11" & x"bf5" => DATA <= x"6000";
            when "11" & x"bf6" => DATA <= x"1d00";
            when "11" & x"bf7" => DATA <= x"03c0";
            when "11" & x"bf8" => DATA <= x"9e00";
            when "11" & x"bf9" => DATA <= x"0100";
            when "11" & x"bfa" => DATA <= x"07c1";
            when "11" & x"bfb" => DATA <= x"e1c0";
            when "11" & x"bfc" => DATA <= x"0540";
            when "11" & x"bfd" => DATA <= x"1080";
            when "11" & x"bfe" => DATA <= x"1404";
            when "11" & x"bff" => DATA <= x"0001";
            when "11" & x"c00" => DATA <= x"0008";
            when "11" & x"c01" => DATA <= x"400a";
            when "11" & x"c02" => DATA <= x"10e0";
            when "11" & x"c03" => DATA <= x"0100";
            when "11" & x"c04" => DATA <= x"0a80";
            when "11" & x"c05" => DATA <= x"011e";
            when "11" & x"c06" => DATA <= x"0140";
            when "11" & x"c07" => DATA <= x"080a";
            when "11" & x"c08" => DATA <= x"0002";
            when "11" & x"c09" => DATA <= x"4803";
            when "11" & x"c0a" => DATA <= x"4020";
            when "11" & x"c0b" => DATA <= x"000a";
            when "11" & x"c0c" => DATA <= x"4802";
            when "11" & x"c0d" => DATA <= x"2e80";
            when "11" & x"c0e" => DATA <= x"1012";
            when "11" & x"c0f" => DATA <= x"0039";
            when "11" & x"c10" => DATA <= x"a004";
            when "11" & x"c11" => DATA <= x"3d00";
            when "11" & x"c12" => DATA <= x"0600";
            when "11" & x"c13" => DATA <= x"0210";
            when "11" & x"c14" => DATA <= x"c000";
            when "11" & x"c15" => DATA <= x"0320";
            when "11" & x"c16" => DATA <= x"020f";
            when "11" & x"c17" => DATA <= x"000c";
            when "11" & x"c18" => DATA <= x"0000";
            when "11" & x"c19" => DATA <= x"2409";
            when "11" & x"c1a" => DATA <= x"0020";
            when "11" & x"c1b" => DATA <= x"5001";
            when "11" & x"c1c" => DATA <= x"97c0";
            when "11" & x"c1d" => DATA <= x"2801";
            when "11" & x"c1e" => DATA <= x"6560";
            when "11" & x"c1f" => DATA <= x"0fc7";
            when "11" & x"c20" => DATA <= x"dbb1";
            when "11" & x"c21" => DATA <= x"f8f8";
            when "11" & x"c22" => DATA <= x"7f57";
            when "11" & x"c23" => DATA <= x"c2fc";
            when "11" & x"c24" => DATA <= x"7f57";
            when "11" & x"c25" => DATA <= x"e3f5";
            when "11" & x"c26" => DATA <= x"ff1f";
            when "11" & x"c27" => DATA <= x"802a";
            when "11" & x"c28" => DATA <= x"5d00";
            when "11" & x"c29" => DATA <= x"b709";
            when "11" & x"c2a" => DATA <= x"0400";
            when "11" & x"c2b" => DATA <= x"2261";
            when "11" & x"c2c" => DATA <= x"0a85";
            when "11" & x"c2d" => DATA <= x"cc00";
            when "11" & x"c2e" => DATA <= x"6338";
            when "11" & x"c2f" => DATA <= x"2b00";
            when "11" & x"c30" => DATA <= x"00ef";
            when "11" & x"c31" => DATA <= x"0600";
            when "11" & x"c32" => DATA <= x"0fa7";
            when "11" & x"c33" => DATA <= x"9452";
            when "11" & x"c34" => DATA <= x"a994";
            when "11" & x"c35" => DATA <= x"e840";
            when "11" & x"c36" => DATA <= x"2290";
            when "11" & x"c37" => DATA <= x"2eaa";
            when "11" & x"c38" => DATA <= x"7f23";
            when "11" & x"c39" => DATA <= x"d3fb";
            when "11" & x"c3a" => DATA <= x"fe9f";
            when "11" & x"c3b" => DATA <= x"df0f";
            when "11" & x"c3c" => DATA <= x"d010";
            when "11" & x"c3d" => DATA <= x"2000";
            when "11" & x"c3e" => DATA <= x"ffa0";
            when "11" & x"c3f" => DATA <= x"077b";
            when "11" & x"c40" => DATA <= x"ff80";
            when "11" & x"c41" => DATA <= x"0074";
            when "11" & x"c42" => DATA <= x"0001";
            when "11" & x"c43" => DATA <= x"0798";
            when "11" & x"c44" => DATA <= x"0013";
            when "11" & x"c45" => DATA <= x"00fc";
            when "11" & x"c46" => DATA <= x"4000";
            when "11" & x"c47" => DATA <= x"00e5";
            when "11" & x"c48" => DATA <= x"f9ff";
            when "11" & x"c49" => DATA <= x"7dbc";
            when "11" & x"c4a" => DATA <= x"0827";
            when "11" & x"c4b" => DATA <= x"0418";
            when "11" & x"c4c" => DATA <= x"edf7";
            when "11" & x"c4d" => DATA <= x"ce20";
            when "11" & x"c4e" => DATA <= x"1000";
            when "11" & x"c4f" => DATA <= x"0400";
            when "11" & x"c50" => DATA <= x"01f0";
            when "11" & x"c51" => DATA <= x"0003";
            when "11" & x"c52" => DATA <= x"beb9";
            when "11" & x"c53" => DATA <= x"fbbe";
            when "11" & x"c54" => DATA <= x"bfc6";
            when "11" & x"c55" => DATA <= x"03e9";
            when "11" & x"c56" => DATA <= x"be1f";
            when "11" & x"c57" => DATA <= x"83f8";
            when "11" & x"c58" => DATA <= x"01fe";
            when "11" & x"c59" => DATA <= x"3f07";
            when "11" & x"c5a" => DATA <= x"801c";
            when "11" & x"c5b" => DATA <= x"1c00";
            when "11" & x"c5c" => DATA <= x"ff30";
            when "11" & x"c5d" => DATA <= x"3c1f";
            when "11" & x"c5e" => DATA <= x"cff7";
            when "11" & x"c5f" => DATA <= x"1109";
            when "11" & x"c60" => DATA <= x"c0c0";
            when "11" & x"c61" => DATA <= x"7057";
            when "11" & x"c62" => DATA <= x"3b3f";
            when "11" & x"c63" => DATA <= x"87c3";
            when "11" & x"c64" => DATA <= x"c174";
            when "11" & x"c65" => DATA <= x"f86c";
            when "11" & x"c66" => DATA <= x"3f44";
            when "11" & x"c67" => DATA <= x"a000";
            when "11" & x"c68" => DATA <= x"2210";
            when "11" & x"c69" => DATA <= x"02a5";
            when "11" & x"c6a" => DATA <= x"a002";
            when "11" & x"c6b" => DATA <= x"252a";
            when "11" & x"c6c" => DATA <= x"37c0";
            when "11" & x"c6d" => DATA <= x"0542";
            when "11" & x"c6e" => DATA <= x"c1fb";
            when "11" & x"c6f" => DATA <= x"bf8f";
            when "11" & x"c70" => DATA <= x"67e7";
            when "11" & x"c71" => DATA <= x"fbf4";
            when "11" & x"c72" => DATA <= x"0008";
            when "11" & x"c73" => DATA <= x"900a";
            when "11" & x"c74" => DATA <= x"ff00";
            when "11" & x"c75" => DATA <= x"0124";
            when "11" & x"c76" => DATA <= x"02bf";
            when "11" & x"c77" => DATA <= x"c001";
            when "11" & x"c78" => DATA <= x"2900";
            when "11" & x"c79" => DATA <= x"aff0";
            when "11" & x"c7a" => DATA <= x"0026";
            when "11" & x"c7b" => DATA <= x"402b";
            when "11" & x"c7c" => DATA <= x"fc00";
            when "11" & x"c7d" => DATA <= x"0490";
            when "11" & x"c7e" => DATA <= x"0aff";
            when "11" & x"c7f" => DATA <= x"0010";
            when "11" & x"c80" => DATA <= x"2402";
            when "11" & x"c81" => DATA <= x"bfc0";
            when "11" & x"c82" => DATA <= x"0a09";
            when "11" & x"c83" => DATA <= x"00af";
            when "11" & x"c84" => DATA <= x"f002";
            when "11" & x"c85" => DATA <= x"4240";
            when "11" & x"c86" => DATA <= x"2bfc";
            when "11" & x"c87" => DATA <= x"2018";
            when "11" & x"c88" => DATA <= x"900a";
            when "11" & x"c89" => DATA <= x"ff10";
            when "11" & x"c8a" => DATA <= x"e805";
            when "11" & x"c8b" => DATA <= x"7fd8";
            when "11" & x"c8c" => DATA <= x"057f";
            when "11" & x"c8d" => DATA <= x"8fc0";
            when "11" & x"c8e" => DATA <= x"2001";
            when "11" & x"c8f" => DATA <= x"fd00";
            when "11" & x"c90" => DATA <= x"57fc";
            when "11" & x"c91" => DATA <= x"8002";
            when "11" & x"c92" => DATA <= x"0015";
            when "11" & x"c93" => DATA <= x"ff20";
            when "11" & x"c94" => DATA <= x"0040";
            when "11" & x"c95" => DATA <= x"057f";
            when "11" & x"c96" => DATA <= x"d805";
            when "11" & x"c97" => DATA <= x"7f84";
            when "11" & x"c98" => DATA <= x"3800";
            when "11" & x"c99" => DATA <= x"2200";
            when "11" & x"c9a" => DATA <= x"affb";
            when "11" & x"c9b" => DATA <= x"00af";
            when "11" & x"c9c" => DATA <= x"fb00";
            when "11" & x"c9d" => DATA <= x"aff0";
            when "11" & x"c9e" => DATA <= x"8680";
            when "11" & x"c9f" => DATA <= x"07df";
            when "11" & x"ca0" => DATA <= x"f600";
            when "11" & x"ca1" => DATA <= x"167f";
            when "11" & x"ca2" => DATA <= x"d803";
            when "11" & x"ca3" => DATA <= x"e1fe";
            when "11" & x"ca4" => DATA <= x"12d0";
            when "11" & x"ca5" => DATA <= x"0aff";
            when "11" & x"ca6" => DATA <= x"b00a";
            when "11" & x"ca7" => DATA <= x"ffb0";
            when "11" & x"ca8" => DATA <= x"07fb";
            when "11" & x"ca9" => DATA <= x"dd01";
            when "11" & x"caa" => DATA <= x"4001";
            when "11" & x"cab" => DATA <= x"25c0";
            when "11" & x"cac" => DATA <= x"02bf";
            when "11" & x"cad" => DATA <= x"ec02";
            when "11" & x"cae" => DATA <= x"bfde";
            when "11" & x"caf" => DATA <= x"1400";
            when "11" & x"cb0" => DATA <= x"8845";
            when "11" & x"cb1" => DATA <= x"022b";
            when "11" & x"cb2" => DATA <= x"fc03";
            when "11" & x"cb3" => DATA <= x"4000";
            when "11" & x"cb4" => DATA <= x"f038";
            when "11" & x"cb5" => DATA <= x"018e";
            when "11" & x"cb6" => DATA <= x"87b0";
            when "11" & x"cb7" => DATA <= x"0aff";
            when "11" & x"cb8" => DATA <= x"b00a";
            when "11" & x"cb9" => DATA <= x"ffb0";
            when "11" & x"cba" => DATA <= x"0aff";
            when "11" & x"cbb" => DATA <= x"b00a";
            when "11" & x"cbc" => DATA <= x"ffb0";
            when "11" & x"cbd" => DATA <= x"07f3";
            when "11" & x"cbe" => DATA <= x"fec0";
            when "11" & x"cbf" => DATA <= x"0fef";
            when "11" & x"cc0" => DATA <= x"f087";
            when "11" & x"cc1" => DATA <= x"0004";
            when "11" & x"cc2" => DATA <= x"000f";
            when "11" & x"cc3" => DATA <= x"c7f8";
            when "11" & x"cc4" => DATA <= x"4380";
            when "11" & x"cc5" => DATA <= x"0220";
            when "11" & x"cc6" => DATA <= x"079b";
            when "11" & x"cc7" => DATA <= x"fec0";
            when "11" & x"cc8" => DATA <= x"1cef";
            when "11" & x"cc9" => DATA <= x"fb00";
            when "11" & x"cca" => DATA <= x"affb";
            when "11" & x"ccb" => DATA <= x"00af";
            when "11" & x"ccc" => DATA <= x"fb00";
            when "11" & x"ccd" => DATA <= x"aff0";
            when "11" & x"cce" => DATA <= x"8700";
            when "11" & x"ccf" => DATA <= x"1800";
            when "11" & x"cd0" => DATA <= x"15ff";
            when "11" & x"cd1" => DATA <= x"2001";
            when "11" & x"cd2" => DATA <= x"f105";
            when "11" & x"cd3" => DATA <= x"7f84";
            when "11" & x"cd4" => DATA <= x"2400";
            when "11" & x"cd5" => DATA <= x"083f";
            when "11" & x"cd6" => DATA <= x"7f8f";
            when "11" & x"cd7" => DATA <= x"b800";
            when "11" & x"cd8" => DATA <= x"fe53";
            when "11" & x"cd9" => DATA <= x"aff0";
            when "11" & x"cda" => DATA <= x"1700";
            when "11" & x"cdb" => DATA <= x"5011";
            when "11" & x"cdc" => DATA <= x"7dff";
            when "11" & x"cdd" => DATA <= x"c001";
            when "11" & x"cde" => DATA <= x"0a00";
            when "11" & x"cdf" => DATA <= x"7e3f";
            when "11" & x"ce0" => DATA <= x"c09c";
            when "11" & x"ce1" => DATA <= x"0020";
            when "11" & x"ce2" => DATA <= x"0057";
            when "11" & x"ce3" => DATA <= x"ff00";
            when "11" & x"ce4" => DATA <= x"1000";
            when "11" & x"ce5" => DATA <= x"4003";
            when "11" & x"ce6" => DATA <= x"fbfe";
            when "11" & x"ce7" => DATA <= x"4000";
            when "11" & x"ce8" => DATA <= x"c00a";
            when "11" & x"ce9" => DATA <= x"ffd0";
            when "11" & x"cea" => DATA <= x"0405";
            when "11" & x"ceb" => DATA <= x"7ff0";
            when "11" & x"cec" => DATA <= x"0006";
            when "11" & x"ced" => DATA <= x"802b";
            when "11" & x"cee" => DATA <= x"fe40";
            when "11" & x"cef" => DATA <= x"0200";
            when "11" & x"cf0" => DATA <= x"0aff";
            when "11" & x"cf1" => DATA <= x"0000";
            when "11" & x"cf2" => DATA <= x"4000";
            when "11" & x"cf3" => DATA <= x"8008";
            when "11" & x"cf4" => DATA <= x"02bf";
            when "11" & x"cf5" => DATA <= x"c000";
            when "11" & x"cf6" => DATA <= x"1a00";
            when "11" & x"cf7" => DATA <= x"0080";
            when "11" & x"cf8" => DATA <= x"2bfe";
            when "11" & x"cf9" => DATA <= x"400b";
            when "11" & x"cfa" => DATA <= x"602a";
            when "11" & x"cfb" => DATA <= x"ff90";
            when "11" & x"cfc" => DATA <= x"0600";
            when "11" & x"cfd" => DATA <= x"02bf";
            when "11" & x"cfe" => DATA <= x"e820";
            when "11" & x"cff" => DATA <= x"00b8";
            when "11" & x"d00" => DATA <= x"0400";
            when "11" & x"d01" => DATA <= x"2bfd";
            when "11" & x"d02" => DATA <= x"fd5f";
            when "11" & x"d03" => DATA <= x"0ff7";
            when "11" & x"d04" => DATA <= x"43f2";
            when "11" & x"d05" => DATA <= x"bfec";
            when "11" & x"d06" => DATA <= x"fd7e";
            when "11" & x"d07" => DATA <= x"3f06";
            when "11" & x"d08" => DATA <= x"3110";
            when "11" & x"d09" => DATA <= x"8c26";
            when "11" & x"d0a" => DATA <= x"2001";
            when "11" & x"d0b" => DATA <= x"8a00";
            when "11" & x"d0c" => DATA <= x"043b";
            when "11" & x"d0d" => DATA <= x"dcf5";
            when "11" & x"d0e" => DATA <= x"ee00";
            when "11" & x"d0f" => DATA <= x"73d0";
            when "11" & x"d10" => DATA <= x"04bc";
            when "11" & x"d11" => DATA <= x"800f";
            when "11" & x"d12" => DATA <= x"2104";
            when "11" & x"d13" => DATA <= x"5555";
            when "11" & x"d14" => DATA <= x"2815";
            when "11" & x"d15" => DATA <= x"4824";
            when "11" & x"d16" => DATA <= x"0ba4";
            when "11" & x"d17" => DATA <= x"8fef";
            when "11" & x"d18" => DATA <= x"e027";
            when "11" & x"d19" => DATA <= x"e1e1";
            when "11" & x"d1a" => DATA <= x"f0c1";
            when "11" & x"d1b" => DATA <= x"6280";
            when "11" & x"d1c" => DATA <= x"0020";
            when "11" & x"d1d" => DATA <= x"07fb";
            when "11" & x"d1e" => DATA <= x"0000";
            when "11" & x"d1f" => DATA <= x"077f";
            when "11" & x"d20" => DATA <= x"bf09";
            when "11" & x"d21" => DATA <= x"0e0a";
            when "11" & x"d22" => DATA <= x"ff7e";
            when "11" & x"d23" => DATA <= x"2000";
            when "11" & x"d24" => DATA <= x"6010";
            when "11" & x"d25" => DATA <= x"06ff";
            when "11" & x"d26" => DATA <= x"bf18";
            when "11" & x"d27" => DATA <= x"000f";
            when "11" & x"d28" => DATA <= x"ff7c";
            when "11" & x"d29" => DATA <= x"5008";
            when "11" & x"d2a" => DATA <= x"475c";
            when "11" & x"d2b" => DATA <= x"4001";
            when "11" & x"d2c" => DATA <= x"0b00";
            when "11" & x"d2d" => DATA <= x"fef7";
            when "11" & x"d2e" => DATA <= x"7808";
            when "11" & x"d2f" => DATA <= x"0002";
            when "11" & x"d30" => DATA <= x"073f";
            when "11" & x"d31" => DATA <= x"a8f9";
            when "11" & x"d32" => DATA <= x"7dc0";
            when "11" & x"d33" => DATA <= x"0fe7";
            when "11" & x"d34" => DATA <= x"f843";
            when "11" & x"d35" => DATA <= x"402b";
            when "11" & x"d36" => DATA <= x"fc3b";
            when "11" & x"d37" => DATA <= x"400e";
            when "11" & x"d38" => DATA <= x"6003";
            when "11" & x"d39" => DATA <= x"81da";
            when "11" & x"d3a" => DATA <= x"ef7a";
            when "11" & x"d3b" => DATA <= x"309c";
            when "11" & x"d3c" => DATA <= x"09f9";
            when "11" & x"d3d" => DATA <= x"1fef";
            when "11" & x"d3e" => DATA <= x"f005";
            when "11" & x"d3f" => DATA <= x"0094";
            when "11" & x"d40" => DATA <= x"0e1d";
            when "11" & x"d41" => DATA <= x"ffc0";
            when "11" & x"d42" => DATA <= x"0a04";
            when "11" & x"d43" => DATA <= x"057f";
            when "11" & x"d44" => DATA <= x"bbdf";
            when "11" & x"d45" => DATA <= x"0c00";
            when "11" & x"d46" => DATA <= x"03e0";
            when "11" & x"d47" => DATA <= x"015f";
            when "11" & x"d48" => DATA <= x"ef77";
            when "11" & x"d49" => DATA <= x"fbbc";
            when "11" & x"d4a" => DATA <= x"147d";
            when "11" & x"d4b" => DATA <= x"003f";
            when "11" & x"d4c" => DATA <= x"d9ef";
            when "11" & x"d4d" => DATA <= x"f6f8";
            when "11" & x"d4e" => DATA <= x"9097";
            when "11" & x"d4f" => DATA <= x"4015";
            when "11" & x"d50" => DATA <= x"fefb";
            when "11" & x"d51" => DATA <= x"7fd0";
            when "11" & x"d52" => DATA <= x"0200";
            when "11" & x"d53" => DATA <= x"015f";
            when "11" & x"d54" => DATA <= x"ef74";
            when "11" & x"d55" => DATA <= x"fd00";
            when "11" & x"d56" => DATA <= x"2bc0";
            when "11" & x"d57" => DATA <= x"0ff7";
            when "11" & x"d58" => DATA <= x"ed7f";
            when "11" & x"d59" => DATA <= x"8802";
            when "11" & x"d5a" => DATA <= x"80f2";
            when "11" & x"d5b" => DATA <= x"057f";
            when "11" & x"d5c" => DATA <= x"bcc0";
            when "11" & x"d5d" => DATA <= x"7201";
            when "11" & x"d5e" => DATA <= x"5fef";
            when "11" & x"d5f" => DATA <= x"d003";
            when "11" & x"d60" => DATA <= x"0110";
            when "11" & x"d61" => DATA <= x"4010";
            when "11" & x"d62" => DATA <= x"57fb";
            when "11" & x"d63" => DATA <= x"ec00";
            when "11" & x"d64" => DATA <= x"7637";
            when "11" & x"d65" => DATA <= x"3fc0";
            when "11" & x"d66" => DATA <= x"15fe";
            when "11" & x"d67" => DATA <= x"fd00";
            when "11" & x"d68" => DATA <= x"1080";
            when "11" & x"d69" => DATA <= x"81f0";
            when "11" & x"d6a" => DATA <= x"03fd";
            when "11" & x"d6b" => DATA <= x"eeff";
            when "11" & x"d6c" => DATA <= x"0003";
            when "11" & x"d6d" => DATA <= x"0034";
            when "11" & x"d6e" => DATA <= x"015f";
            when "11" & x"d6f" => DATA <= x"efee";
            when "11" & x"d70" => DATA <= x"0052";
            when "11" & x"d71" => DATA <= x"005f";
            when "11" & x"d72" => DATA <= x"e7f7";
            when "11" & x"d73" => DATA <= x"cb02";
            when "11" & x"d74" => DATA <= x"801f";
            when "11" & x"d75" => DATA <= x"c00a";
            when "11" & x"d76" => DATA <= x"ff7f";
            when "11" & x"d77" => DATA <= x"0dd6";
            when "11" & x"d78" => DATA <= x"0040";
            when "11" & x"d79" => DATA <= x"1842";
            when "11" & x"d7a" => DATA <= x"bfcf";
            when "11" & x"d7b" => DATA <= x"c007";
            when "11" & x"d7c" => DATA <= x"9182";
            when "11" & x"d7d" => DATA <= x"803b";
            when "11" & x"d7e" => DATA <= x"fc02";
            when "11" & x"d7f" => DATA <= x"6751";
            when "11" & x"d80" => DATA <= x"b700";
            when "11" & x"d81" => DATA <= x"15fe";
            when "11" & x"d82" => DATA <= x"7f02";
            when "11" & x"d83" => DATA <= x"09eb";
            when "11" & x"d84" => DATA <= x"fc01";
            when "11" & x"d85" => DATA <= x"dfe0";
            when "11" & x"d86" => DATA <= x"0109";
            when "11" & x"d87" => DATA <= x"fc0e";
            when "11" & x"d88" => DATA <= x"007f";
            when "11" & x"d89" => DATA <= x"bf57";
            when "11" & x"d8a" => DATA <= x"e000";
            when "11" & x"d8b" => DATA <= x"0afc";
            when "11" & x"d8c" => DATA <= x"0001";
            when "11" & x"d8d" => DATA <= x"eff7";
            when "11" & x"d8e" => DATA <= x"c001";
            when "11" & x"d8f" => DATA <= x"fefa";
            when "11" & x"d90" => DATA <= x"003f";
            when "11" & x"d91" => DATA <= x"dbef";
            when "11" & x"d92" => DATA <= x"e018";
            when "11" & x"d93" => DATA <= x"006e";
            when "11" & x"d94" => DATA <= x"ff00";
            when "11" & x"d95" => DATA <= x"57fa";
            when "11" & x"d96" => DATA <= x"fcd8";
            when "11" & x"d97" => DATA <= x"d409";
            when "11" & x"d98" => DATA <= x"5005";
            when "11" & x"d99" => DATA <= x"7fb7";
            when "11" & x"d9a" => DATA <= x"df2b";
            when "11" & x"d9b" => DATA <= x"f495";
            when "11" & x"d9c" => DATA <= x"0057";
            when "11" & x"d9d" => DATA <= x"f9fd";
            when "11" & x"d9e" => DATA <= x"fefb";
            when "11" & x"d9f" => DATA <= x"2e39";
            when "11" & x"da0" => DATA <= x"0015";
            when "11" & x"da1" => DATA <= x"fedf";
            when "11" & x"da2" => DATA <= x"7f8b";
            when "11" & x"da3" => DATA <= x"c84f";
            when "11" & x"da4" => DATA <= x"f003";
            when "11" & x"da5" => DATA <= x"fcff";
            when "11" & x"da6" => DATA <= x"5fe4";
            when "11" & x"da7" => DATA <= x"2048";
            when "11" & x"da8" => DATA <= x"0c01";
            when "11" & x"da9" => DATA <= x"5fee";
            when "11" & x"daa" => DATA <= x"e7fc";
            when "11" & x"dab" => DATA <= x"e07f";
            when "11" & x"dac" => DATA <= x"fcff";
            when "11" & x"dad" => DATA <= x"f43b";
            when "11" & x"dae" => DATA <= x"1e61";
            when "11" & x"daf" => DATA <= x"ffff";
            when "11" & x"db0" => DATA <= x"bffb";
            when "11" & x"db1" => DATA <= x"cfb8";
            when "11" & x"db2" => DATA <= x"ebfc";
            when "11" & x"db3" => DATA <= x"6bff";
            when "11" & x"db4" => DATA <= x"e007";
            when "11" & x"db5" => DATA <= x"38ff";
            when "11" & x"db6" => DATA <= x"7fc0";
            when "11" & x"db7" => DATA <= x"0782";
            when "11" & x"db8" => DATA <= x"057f";
            when "11" & x"db9" => DATA <= x"bdeb";
            when "11" & x"dba" => DATA <= x"fc42";
            when "11" & x"dbb" => DATA <= x"fe00";
            when "11" & x"dbc" => DATA <= x"57fb";
            when "11" & x"dbd" => DATA <= x"eebf";
            when "11" & x"dbe" => DATA <= x"d483";
            when "11" & x"dbf" => DATA <= x"f003";
            when "11" & x"dc0" => DATA <= x"fdcf";
            when "11" & x"dc1" => DATA <= x"dfe0";
            when "11" & x"dc2" => DATA <= x"b7f8";
            when "11" & x"dc3" => DATA <= x"12bf";
            when "11" & x"dc4" => DATA <= x"dfb5";
            when "11" & x"dc5" => DATA <= x"fe00";
            when "11" & x"dc6" => DATA <= x"6780";
            when "11" & x"dc7" => DATA <= x"2bfd";
            when "11" & x"dc8" => DATA <= x"f75f";
            when "11" & x"dc9" => DATA <= x"e007";
            when "11" & x"dca" => DATA <= x"f803";
            when "11" & x"dcb" => DATA <= x"7fc0";
            when "11" & x"dcc" => DATA <= x"0270";
            when "11" & x"dcd" => DATA <= x"057f";
            when "11" & x"dce" => DATA <= x"bf7b";
            when "11" & x"dcf" => DATA <= x"fdce";
            when "11" & x"dd0" => DATA <= x"00af";
            when "11" & x"dd1" => DATA <= x"f7f5";
            when "11" & x"dd2" => DATA <= x"7faf";
            when "11" & x"dd3" => DATA <= x"d3c1";
            when "11" & x"dd4" => DATA <= x"0aff";
            when "11" & x"dd5" => DATA <= x"7ecf";
            when "11" & x"dd6" => DATA <= x"f802";
            when "11" & x"dd7" => DATA <= x"bfdf";
            when "11" & x"dd8" => DATA <= x"ddfe";
            when "11" & x"dd9" => DATA <= x"0f00";
            when "11" & x"dda" => DATA <= x"3fdf";
            when "11" & x"ddb" => DATA <= x"27fe";
            when "11" & x"ddc" => DATA <= x"ff20";
            when "11" & x"ddd" => DATA <= x"382f";
            when "11" & x"dde" => DATA <= x"fdf0";
            when "11" & x"ddf" => DATA <= x"f0ff";
            when "11" & x"de0" => DATA <= x"ffff";
            when "11" & x"de1" => DATA <= x"fff1";
            when "11" & x"de2" => DATA <= x"fafe";
            when "11" & x"de3" => DATA <= x"ffcb";
            when "11" & x"de4" => DATA <= x"200b";
            when "11" & x"de5" => DATA <= x"ff01";
            when "11" & x"de6" => DATA <= x"803b";
            when "11" & x"de7" => DATA <= x"fc01";
            when "11" & x"de8" => DATA <= x"5fef";
            when "11" & x"de9" => DATA <= x"c707";
            when "11" & x"dea" => DATA <= x"7f80";
            when "11" & x"deb" => DATA <= x"2bfc";
            when "11" & x"dec" => DATA <= x"fb3f";
            when "11" & x"ded" => DATA <= x"e01a";
            when "11" & x"dee" => DATA <= x"ff01";
            when "11" & x"def" => DATA <= x"1feb";
            when "11" & x"df0" => DATA <= x"fdf6";
            when "11" & x"df1" => DATA <= x"04af";
            when "11" & x"df2" => DATA <= x"fa00";
            when "11" & x"df3" => DATA <= x"aff6";
            when "11" & x"df4" => DATA <= x"6831";
            when "11" & x"df5" => DATA <= x"fefe";
            when "11" & x"df6" => DATA <= x"1077";
            when "11" & x"df7" => DATA <= x"fbdc";
            when "11" & x"df8" => DATA <= x"015f";
            when "11" & x"df9" => DATA <= x"e7d9";
            when "11" & x"dfa" => DATA <= x"ff00";
            when "11" & x"dfb" => DATA <= x"57fb";
            when "11" & x"dfc" => DATA <= x"91c3";
            when "11" & x"dfd" => DATA <= x"dfe0";
            when "11" & x"dfe" => DATA <= x"0eff";
            when "11" & x"dff" => DATA <= x"03f7";
            when "11" & x"e00" => DATA <= x"f902";
            when "11" & x"e01" => DATA <= x"afc7";
            when "11" & x"e02" => DATA <= x"f3ff";
            when "11" & x"e03" => DATA <= x"c00f";
            when "11" & x"e04" => DATA <= x"6787";
            when "11" & x"e05" => DATA <= x"7fa0";
            when "11" & x"e06" => DATA <= x"1f00";
            when "11" & x"e07" => DATA <= x"04b9";
            when "11" & x"e08" => DATA <= x"57bf";
            when "11" & x"e09" => DATA <= x"c000";
            when "11" & x"e0a" => DATA <= x"3000";
            when "11" & x"e0b" => DATA <= x"183c";
            when "11" & x"e0c" => DATA <= x"ff7b";
            when "11" & x"e0d" => DATA <= x"bf40";
            when "11" & x"e0e" => DATA <= x"0a94";
            when "11" & x"e0f" => DATA <= x"6a01";
            when "11" & x"e10" => DATA <= x"047f";
            when "11" & x"e11" => DATA <= x"7fbd";
            when "11" & x"e12" => DATA <= x"80da";
            when "11" & x"e13" => DATA <= x"fe7e";
            when "11" & x"e14" => DATA <= x"7dd0";
            when "11" & x"e15" => DATA <= x"0180";
            when "11" & x"e16" => DATA <= x"0840";
            when "11" & x"e17" => DATA <= x"0200";
            when "11" & x"e18" => DATA <= x"002f";
            when "11" & x"e19" => DATA <= x"f025";
            when "11" & x"e1a" => DATA <= x"0001";
            when "11" & x"e1b" => DATA <= x"2801";
            when "11" & x"e1c" => DATA <= x"803f";
            when "11" & x"e1d" => DATA <= x"a800";
            when "11" & x"e1e" => DATA <= x"0200";
            when "11" & x"e1f" => DATA <= x"0040";
            when "11" & x"e20" => DATA <= x"2110";
            when "11" & x"e21" => DATA <= x"00e0";
            when "11" & x"e22" => DATA <= x"f9ff";
            when "11" & x"e23" => DATA <= x"afe7";
            when "11" & x"e24" => DATA <= x"0000";
            when "11" & x"e25" => DATA <= x"c003";
            when "11" & x"e26" => DATA <= x"3df7";
            when "11" & x"e27" => DATA <= x"f9c4";
            when "11" & x"e28" => DATA <= x"c200";
            when "11" & x"e29" => DATA <= x"0080";
            when "11" & x"e2a" => DATA <= x"3807";
            when "11" & x"e2b" => DATA <= x"c003";
            when "11" & x"e2c" => DATA <= x"8efb";
            when "11" & x"e2d" => DATA <= x"ff77";
            when "11" & x"e2e" => DATA <= x"afaa";
            when "11" & x"e2f" => DATA <= x"ff8f";
            when "11" & x"e30" => DATA <= x"80c3";
            when "11" & x"e31" => DATA <= x"27f8";
            when "11" & x"e32" => DATA <= x"7c4e";
            when "11" & x"e33" => DATA <= x"0060";
            when "11" & x"e34" => DATA <= x"7005";
            when "11" & x"e35" => DATA <= x"3e3e";
            when "11" & x"e36" => DATA <= x"2bfc";
            when "11" & x"e37" => DATA <= x"0150";
            when "11" & x"e38" => DATA <= x"0c07";
            when "11" & x"e39" => DATA <= x"038d";
            when "11" & x"e3a" => DATA <= x"cedf";
            when "11" & x"e3b" => DATA <= x"6391";
            when "11" & x"e3c" => DATA <= x"dfe1";
            when "11" & x"e3d" => DATA <= x"f0ba";
            when "11" & x"e3e" => DATA <= x"7f87";
            when "11" & x"e3f" => DATA <= x"c1cf";
            when "11" & x"e40" => DATA <= x"f780";
            when "11" & x"e41" => DATA <= x"0807";
            when "11" & x"e42" => DATA <= x"4054";
            when "11" & x"e43" => DATA <= x"0027";
            when "11" & x"e44" => DATA <= x"0080";
            when "11" & x"e45" => DATA <= x"0020";
            when "11" & x"e46" => DATA <= x"0008";
            when "11" & x"e47" => DATA <= x"0280";
            when "11" & x"e48" => DATA <= x"4015";
            when "11" & x"e49" => DATA <= x"fc1e";
            when "11" & x"e4a" => DATA <= x"a06a";
            when "11" & x"e4b" => DATA <= x"80a0";
            when "11" & x"e4c" => DATA <= x"03c0";
            when "11" & x"e4d" => DATA <= x"e0f8";
            when "11" & x"e4e" => DATA <= x"7e3f";
            when "11" & x"e4f" => DATA <= x"bfd0";
            when "11" & x"e50" => DATA <= x"004d";
            when "11" & x"e51" => DATA <= x"001b";
            when "11" & x"e52" => DATA <= x"8000";
            when "11" & x"e53" => DATA <= x"5a00";
            when "11" & x"e54" => DATA <= x"1200";
            when "11" & x"e55" => DATA <= x"3003";
            when "11" & x"e56" => DATA <= x"e030";
            when "11" & x"e57" => DATA <= x"0b05";
            when "11" & x"e58" => DATA <= x"e070";
            when "11" & x"e59" => DATA <= x"0007";
            when "11" & x"e5a" => DATA <= x"e87b";
            when "11" & x"e5b" => DATA <= x"87c0";
            when "11" & x"e5c" => DATA <= x"1480";
            when "11" & x"e5d" => DATA <= x"4800";
            when "11" & x"e5e" => DATA <= x"7201";
            when "11" & x"e5f" => DATA <= x"2001";
            when "11" & x"e60" => DATA <= x"b01c";
            when "11" & x"e61" => DATA <= x"003f";
            when "11" & x"e62" => DATA <= x"0780";
            when "11" & x"e63" => DATA <= x"d02c";
            when "11" & x"e64" => DATA <= x"1ae0";
            when "11" & x"e65" => DATA <= x"a00d";
            when "11" & x"e66" => DATA <= x"1f7f";
            when "11" & x"e67" => DATA <= x"8828";
            when "11" & x"e68" => DATA <= x"0101";
            when "11" & x"e69" => DATA <= x"c008";
            when "11" & x"e6a" => DATA <= x"da00";
            when "11" & x"e6b" => DATA <= x"9c02";
            when "11" & x"e6c" => DATA <= x"00f8";
            when "11" & x"e6d" => DATA <= x"00f0";
            when "11" & x"e6e" => DATA <= x"61a0";
            when "11" & x"e6f" => DATA <= x"180e";
            when "11" & x"e70" => DATA <= x"0780";
            when "11" & x"e71" => DATA <= x"4001";
            when "11" & x"e72" => DATA <= x"60e0";
            when "11" & x"e73" => DATA <= x"0e10";
            when "11" & x"e74" => DATA <= x"0048";
            when "11" & x"e75" => DATA <= x"8001";
            when "11" & x"e76" => DATA <= x"c060";
            when "11" & x"e77" => DATA <= x"a203";
            when "11" & x"e78" => DATA <= x"0082";
            when "11" & x"e79" => DATA <= x"8002";
            when "11" & x"e7a" => DATA <= x"0f0a";
            when "11" & x"e7b" => DATA <= x"e0ef";
            when "11" & x"e7c" => DATA <= x"0001";
            when "11" & x"e7d" => DATA <= x"000e";
            when "11" & x"e7e" => DATA <= x"47e0";
            when "11" & x"e7f" => DATA <= x"73f8";
            when "11" & x"e80" => DATA <= x"22c0";
            when "11" & x"e81" => DATA <= x"0c60";
            when "11" & x"e82" => DATA <= x"0009";
            when "11" & x"e83" => DATA <= x"c29c";
            when "11" & x"e84" => DATA <= x"6bc0";
            when "11" & x"e85" => DATA <= x"7e00";
            when "11" & x"e86" => DATA <= x"7c3c";
            when "11" & x"e87" => DATA <= x"2b81";
            when "11" & x"e88" => DATA <= x"e0e0";
            when "11" & x"e89" => DATA <= x"a00d";
            when "11" & x"e8a" => DATA <= x"0300";
            when "11" & x"e8b" => DATA <= x"8000";
            when "11" & x"e8c" => DATA <= x"8440";
            when "11" & x"e8d" => DATA <= x"2002";
            when "11" & x"e8e" => DATA <= x"4100";
            when "11" & x"e8f" => DATA <= x"0b8e";
            when "11" & x"e90" => DATA <= x"181c";
            when "11" & x"e91" => DATA <= x"1e28";
            when "11" & x"e92" => DATA <= x"000e";
            when "11" & x"e93" => DATA <= x"fc7c";
            when "11" & x"e94" => DATA <= x"7783";
            when "11" & x"e95" => DATA <= x"8280";
            when "11" & x"e96" => DATA <= x"3405";
            when "11" & x"e97" => DATA <= x"bf5c";
            when "11" & x"e98" => DATA <= x"460a";
            when "11" & x"e99" => DATA <= x"e270";
            when "11" & x"e9a" => DATA <= x"3000";
            when "11" & x"e9b" => DATA <= x"15fe";
            when "11" & x"e9c" => DATA <= x"f870";
            when "11" & x"e9d" => DATA <= x"3010";
            when "11" & x"e9e" => DATA <= x"2830";
            when "11" & x"e9f" => DATA <= x"17c3";
            when "11" & x"ea0" => DATA <= x"a03f";
            when "11" & x"ea1" => DATA <= x"fdff";
            when "11" & x"ea2" => DATA <= x"fc60";
            when "11" & x"ea3" => DATA <= x"3aff";
            when "11" & x"ea4" => DATA <= x"70a0";
            when "11" & x"ea5" => DATA <= x"4060";
            when "11" & x"ea6" => DATA <= x"7078";
            when "11" & x"ea7" => DATA <= x"188e";
            when "11" & x"ea8" => DATA <= x"0723";
            when "11" & x"ea9" => DATA <= x"81e9";
            when "11" & x"eaa" => DATA <= x"1c8c";
            when "11" & x"eab" => DATA <= x"40a0";
            when "11" & x"eac" => DATA <= x"0010";
            when "11" & x"ead" => DATA <= x"0005";
            when "11" & x"eae" => DATA <= x"4000";
            when "11" & x"eaf" => DATA <= x"2001";
            when "11" & x"eb0" => DATA <= x"fd8e";
            when "11" & x"eb1" => DATA <= x"071b";
            when "11" & x"eb2" => DATA <= x"83c7";
            when "11" & x"eb3" => DATA <= x"e40a";
            when "11" & x"eb4" => DATA <= x"000f";
            when "11" & x"eb5" => DATA <= x"87a8";
            when "11" & x"eb6" => DATA <= x"7030";
            when "11" & x"eb7" => DATA <= x"f030";
            when "11" & x"eb8" => DATA <= x"5800";
            when "11" & x"eb9" => DATA <= x"2d20";
            when "11" & x"eba" => DATA <= x"0440";
            when "11" & x"ebb" => DATA <= x"5425";
            when "11" & x"ebc" => DATA <= x"403f";
            when "11" & x"ebd" => DATA <= x"400e";
            when "11" & x"ebe" => DATA <= x"070d";
            when "11" & x"ebf" => DATA <= x"0183";
            when "11" & x"ec0" => DATA <= x"e8fc";
            when "11" & x"ec1" => DATA <= x"11c1";
            when "11" & x"ec2" => DATA <= x"e0e0";
            when "11" & x"ec3" => DATA <= x"6020";
            when "11" & x"ec4" => DATA <= x"0030";
            when "11" & x"ec5" => DATA <= x"082c";
            when "11" & x"ec6" => DATA <= x"000b";
            when "11" & x"ec7" => DATA <= x"4080";
            when "11" & x"ec8" => DATA <= x"c168";
            when "11" & x"ec9" => DATA <= x"0060";
            when "11" & x"eca" => DATA <= x"0008";
            when "11" & x"ecb" => DATA <= x"1d81";
            when "11" & x"ecc" => DATA <= x"4001";
            when "11" & x"ecd" => DATA <= x"f7c3";
            when "11" & x"ece" => DATA <= x"0002";
            when "11" & x"ecf" => DATA <= x"070f";
            when "11" & x"ed0" => DATA <= x"f004";
            when "11" & x"ed1" => DATA <= x"8381";
            when "11" & x"ed2" => DATA <= x"1f8f";
            when "11" & x"ed3" => DATA <= x"8080";
            when "11" & x"ed4" => DATA <= x"0284";
            when "11" & x"ed5" => DATA <= x"2800";
            when "11" & x"ed6" => DATA <= x"04ff";
            when "11" & x"ed7" => DATA <= x"0030";
            when "11" & x"ed8" => DATA <= x"c0e0";
            when "11" & x"ed9" => DATA <= x"f3ff";
            when "11" & x"eda" => DATA <= x"7f80";
            when "11" & x"edb" => DATA <= x"07ef";
            when "11" & x"edc" => DATA <= x"c783";
            when "11" & x"edd" => DATA <= x"8002";
            when "11" & x"ede" => DATA <= x"037f";
            when "11" & x"edf" => DATA <= x"8018";
            when "11" & x"ee0" => DATA <= x"1dff";
            when "11" & x"ee1" => DATA <= x"580f";
            when "11" & x"ee2" => DATA <= x"f003";
            when "11" & x"ee3" => DATA <= x"c102";
            when "11" & x"ee4" => DATA <= x"0307";
            when "11" & x"ee5" => DATA <= x"9fdf";
            when "11" & x"ee6" => DATA <= x"e7f4";
            when "11" & x"ee7" => DATA <= x"001c";
            when "11" & x"ee8" => DATA <= x"1e0e";
            when "11" & x"ee9" => DATA <= x"4670";
            when "11" & x"eea" => DATA <= x"0028";
            when "11" & x"eeb" => DATA <= x"0080";
            when "11" & x"eec" => DATA <= x"9000";
            when "11" & x"eed" => DATA <= x"8001";
            when "11" & x"eee" => DATA <= x"301f";
            when "11" & x"eef" => DATA <= x"1fbf";
            when "11" & x"ef0" => DATA <= x"df00";
            when "11" & x"ef1" => DATA <= x"0603";
            when "11" & x"ef2" => DATA <= x"f1fe";
            when "11" & x"ef3" => DATA <= x"f060";
            when "11" & x"ef4" => DATA <= x"2001";
            when "11" & x"ef5" => DATA <= x"e1c0";
            when "11" & x"ef6" => DATA <= x"0004";
            when "11" & x"ef7" => DATA <= x"23c0";
            when "11" & x"ef8" => DATA <= x"2006";
            when "11" & x"ef9" => DATA <= x"e022";
            when "11" & x"efa" => DATA <= x"8324";
            when "11" & x"efb" => DATA <= x"0147";
            when "11" & x"efc" => DATA <= x"5800";
            when "11" & x"efd" => DATA <= x"2607";
            when "11" & x"efe" => DATA <= x"613f";
            when "11" & x"eff" => DATA <= x"8020";
            when "11" & x"f00" => DATA <= x"f7c2";
            when "11" & x"f01" => DATA <= x"0002";
            when "11" & x"f02" => DATA <= x"1f3f";
            when "11" & x"f03" => DATA <= x"87c0";
            when "11" & x"f04" => DATA <= x"4000";
            when "11" & x"f05" => DATA <= x"39fc";
            when "11" & x"f06" => DATA <= x"fc78";
            when "11" & x"f07" => DATA <= x"a005";
            when "11" & x"f08" => DATA <= x"0043";
            when "11" & x"f09" => DATA <= x"8002";
            when "11" & x"f0a" => DATA <= x"1c00";
            when "11" & x"f0b" => DATA <= x"0500";
            when "11" & x"f0c" => DATA <= x"7605";
            when "11" & x"f0d" => DATA <= x"0002";
            when "11" & x"f0e" => DATA <= x"000c";
            when "11" & x"f0f" => DATA <= x"4078";
            when "11" & x"f10" => DATA <= x"fdfe";
            when "11" & x"f11" => DATA <= x"fc00";
            when "11" & x"f12" => DATA <= x"1c1f";
            when "11" & x"f13" => DATA <= x"cff7";
            when "11" & x"f14" => DATA <= x"8300";
            when "11" & x"f15" => DATA <= x"021f";
            when "11" & x"f16" => DATA <= x"1f50";
            when "11" & x"f17" => DATA <= x"0022";
            when "11" & x"f18" => DATA <= x"4010";
            when "11" & x"f19" => DATA <= x"000a";
            when "11" & x"f1a" => DATA <= x"0690";
            when "11" & x"f1b" => DATA <= x"0285";
            when "11" & x"f1c" => DATA <= x"0020";
            when "11" & x"f1d" => DATA <= x"4006";
            when "11" & x"f1e" => DATA <= x"170b";
            when "11" & x"f1f" => DATA <= x"c5ff";
            when "11" & x"f20" => DATA <= x"400f";
            when "11" & x"f21" => DATA <= x"f600";
            when "11" & x"f22" => DATA <= x"007e";
            when "11" & x"f23" => DATA <= x"ff03";
            when "11" & x"f24" => DATA <= x"d000";
            when "11" & x"f25" => DATA <= x"0c3e";
            when "11" & x"f26" => DATA <= x"fe70";
            when "11" & x"f27" => DATA <= x"0040";
            when "11" & x"f28" => DATA <= x"0403";
            when "11" & x"f29" => DATA <= x"83c1";
            when "11" & x"f2a" => DATA <= x"fd5f";
            when "11" & x"f2b" => DATA <= x"f501";
            when "11" & x"f2c" => DATA <= x"ffff";
            when "11" & x"f2d" => DATA <= x"ff5f";
            when "11" & x"f2e" => DATA <= x"fee2";
            when "11" & x"f2f" => DATA <= x"710e";
            when "11" & x"f30" => DATA <= x"7804";
            when "11" & x"f31" => DATA <= x"f7d7";
            when "11" & x"f32" => DATA <= x"fd00";
            when "11" & x"f33" => DATA <= x"2f1f";
            when "11" & x"f34" => DATA <= x"d3fe";
            when "11" & x"f35" => DATA <= x"0060";
            when "11" & x"f36" => DATA <= x"5ff8";
            when "11" & x"f37" => DATA <= x"03ff";
            when "11" & x"f38" => DATA <= x"c01f";
            when "11" & x"f39" => DATA <= x"fe00";
            when "11" & x"f3a" => DATA <= x"0fdf";
            when "11" & x"f3b" => DATA <= x"fd00";
            when "11" & x"f3c" => DATA <= x"36f7";
            when "11" & x"f3d" => DATA <= x"fe80";
            when "11" & x"f3e" => DATA <= x"0042";
            when "11" & x"f3f" => DATA <= x"11ff";
            when "11" & x"f40" => DATA <= x"7fd0";
            when "11" & x"f41" => DATA <= x"03c1";
            when "11" & x"f42" => DATA <= x"f0fe";
            when "11" & x"f43" => DATA <= x"effa";
            when "11" & x"f44" => DATA <= x"00bf";
            when "11" & x"f45" => DATA <= x"fa00";
            when "11" & x"f46" => DATA <= x"bffa";
            when "11" & x"f47" => DATA <= x"0002";
            when "11" & x"f48" => DATA <= x"9ce7";
            when "11" & x"f49" => DATA <= x"fe80";
            when "11" & x"f4a" => DATA <= x"1f0f";
            when "11" & x"f4b" => DATA <= x"e9ff";
            when "11" & x"f4c" => DATA <= x"003f";
            when "11" & x"f4d" => DATA <= x"2ffc";
            when "11" & x"f4e" => DATA <= x"0001";
            when "11" & x"f4f" => DATA <= x"5ad7";
            when "11" & x"f50" => DATA <= x"f9fc";
            when "11" & x"f51" => DATA <= x"7ec7";
            when "11" & x"f52" => DATA <= x"a000";
            when "11" & x"f53" => DATA <= x"1004";
            when "11" & x"f54" => DATA <= x"0084";
            when "11" & x"f55" => DATA <= x"61bc";
            when "11" & x"f56" => DATA <= x"4008";
            when "11" & x"f57" => DATA <= x"07c3";
            when "11" & x"f58" => DATA <= x"fa7f";
            when "11" & x"f59" => DATA <= x"c01f";
            when "11" & x"f5a" => DATA <= x"fe00";
            when "11" & x"f5b" => DATA <= x"07df";
            when "11" & x"f5c" => DATA <= x"fd00";
            when "11" & x"f5d" => DATA <= x"07db";
            when "11" & x"f5e" => DATA <= x"f3ff";
            when "11" & x"f5f" => DATA <= x"400f";
            when "11" & x"f60" => DATA <= x"07cc";
            when "11" & x"f61" => DATA <= x"ffd0";
            when "11" & x"f62" => DATA <= x"01ff";
            when "11" & x"f63" => DATA <= x"7fc0";
            when "11" & x"f64" => DATA <= x"0ff3";
            when "11" & x"f65" => DATA <= x"6eff";
            when "11" & x"f66" => DATA <= x"8000";
            when "11" & x"f67" => DATA <= x"20d4";
            when "11" & x"f68" => DATA <= x"7b3f";
            when "11" & x"f69" => DATA <= x"bfe8";
            when "11" & x"f6a" => DATA <= x"01e0";
            when "11" & x"f6b" => DATA <= x"f17d";
            when "11" & x"f6c" => DATA <= x"bf6b";
            when "11" & x"f6d" => DATA <= x"fe80";
            when "11" & x"f6e" => DATA <= x"2ffc";
            when "11" & x"f6f" => DATA <= x"00f0";
            when "11" & x"f70" => DATA <= x"bff0";
            when "11" & x"f71" => DATA <= x"007c";
            when "11" & x"f72" => DATA <= x"7fcf";
            when "11" & x"f73" => DATA <= x"f5ff";
            when "11" & x"f74" => DATA <= x"400e";
            when "11" & x"f75" => DATA <= x"0733";
            when "11" & x"f76" => DATA <= x"1ddf";
            when "11" & x"f77" => DATA <= x"5ff4";
            when "11" & x"f78" => DATA <= x"005f";
            when "11" & x"f79" => DATA <= x"dffa";
            when "11" & x"f7a" => DATA <= x"002d";
            when "11" & x"f7b" => DATA <= x"6ff8";
            when "11" & x"f7c" => DATA <= x"001f";
            when "11" & x"f7d" => DATA <= x"47e7";
            when "11" & x"f7e" => DATA <= x"feff";
            when "11" & x"f7f" => DATA <= x"a007";
            when "11" & x"f80" => DATA <= x"038a";
            when "11" & x"f81" => DATA <= x"bdeb";
            when "11" & x"f82" => DATA <= x"fe80";
            when "11" & x"f83" => DATA <= x"2ffc";
            when "11" & x"f84" => DATA <= x"00e0";
            when "11" & x"f85" => DATA <= x"77ef";
            when "11" & x"f86" => DATA <= x"f802";
            when "11" & x"f87" => DATA <= x"80c0";
            when "11" & x"f88" => DATA <= x"2311";
            when "11" & x"f89" => DATA <= x"99cc";
            when "11" & x"f8a" => DATA <= x"ff40";
            when "11" & x"f8b" => DATA <= x"0efa";
            when "11" & x"f8c" => DATA <= x"feef";
            when "11" & x"f8d" => DATA <= x"fa00";
            when "11" & x"f8e" => DATA <= x"bff0";
            when "11" & x"f8f" => DATA <= x"03f9";
            when "11" & x"f90" => DATA <= x"dfbf";
            when "11" & x"f91" => DATA <= x"f401";
            when "11" & x"f92" => DATA <= x"4063";
            when "11" & x"f93" => DATA <= x"31da";
            when "11" & x"f94" => DATA <= x"edff";
            when "11" & x"f95" => DATA <= x"400e";
            when "11" & x"f96" => DATA <= x"e7e3";
            when "11" & x"f97" => DATA <= x"fbbf";
            when "11" & x"f98" => DATA <= x"c008";
            when "11" & x"f99" => DATA <= x"07ae";
            when "11" & x"f9a" => DATA <= x"ff80";
            when "11" & x"f9b" => DATA <= x"1fe7";
            when "11" & x"f9c" => DATA <= x"fa3f";
            when "11" & x"f9d" => DATA <= x"0f8f";
            when "11" & x"f9e" => DATA <= x"c3f4";
            when "11" & x"f9f" => DATA <= x"00f0";
            when "11" & x"fa0" => DATA <= x"9e06";
            when "11" & x"fa1" => DATA <= x"1d00";
            when "11" & x"fa2" => DATA <= x"5ff8";
            when "11" & x"fa3" => DATA <= x"01f1";
            when "11" & x"fa4" => DATA <= x"7fe0";
            when "11" & x"fa5" => DATA <= x"07ff";
            when "11" & x"fa6" => DATA <= x"1ff0";
            when "11" & x"fa7" => DATA <= x"fd00";
            when "11" & x"fa8" => DATA <= x"1c3b";
            when "11" & x"fa9" => DATA <= x"c1e2";
            when "11" & x"faa" => DATA <= x"f0a0";
            when "11" & x"fab" => DATA <= x"03de";
            when "11" & x"fac" => DATA <= x"ff80";
            when "11" & x"fad" => DATA <= x"1fef";
            when "11" & x"fae" => DATA <= x"bdff";
            when "11" & x"faf" => DATA <= x"003f";
            when "11" & x"fb0" => DATA <= x"c1f4";
            when "11" & x"fb1" => DATA <= x"3fc1";
            when "11" & x"fb2" => DATA <= x"e000";
            when "11" & x"fb3" => DATA <= x"0d7c";
            when "11" & x"fb4" => DATA <= x"7783";
            when "11" & x"fb5" => DATA <= x"8680";
            when "11" & x"fb6" => DATA <= x"2ffc";
            when "11" & x"fb7" => DATA <= x"00fe";
            when "11" & x"fb8" => DATA <= x"bff0";
            when "11" & x"fb9" => DATA <= x"03fc";
            when "11" & x"fba" => DATA <= x"0740";
            when "11" & x"fbb" => DATA <= x"fc1e";
            when "11" & x"fbc" => DATA <= x"0001";
            when "11" & x"fbd" => DATA <= x"bfeb";
            when "11" & x"fbe" => DATA <= x"f9f8";
            when "11" & x"fbf" => DATA <= x"f878";
            when "11" & x"fc0" => DATA <= x"5005";
            when "11" & x"fc1" => DATA <= x"ff80";
            when "11" & x"fc2" => DATA <= x"1fec";
            when "11" & x"fc3" => DATA <= x"040d";
            when "11" & x"fc4" => DATA <= x"01d0";
            when "11" & x"fc5" => DATA <= x"3800";
            when "11" & x"fc6" => DATA <= x"03df";
            when "11" & x"fc7" => DATA <= x"efe7";
            when "11" & x"fc8" => DATA <= x"e3e0";
            when "11" & x"fc9" => DATA <= x"0080";
            when "11" & x"fca" => DATA <= x"bff0";
            when "11" & x"fcb" => DATA <= x"03fe";
            when "11" & x"fcc" => DATA <= x"8fcf";
            when "11" & x"fcd" => DATA <= x"fdfe";
            when "11" & x"fce" => DATA <= x"007f";
            when "11" & x"fcf" => DATA <= x"be1e";
            when "11" & x"fd0" => DATA <= x"0e06";
            when "11" & x"fd1" => DATA <= x"0200";
            when "11" & x"fd2" => DATA <= x"0340";
            when "11" & x"fd3" => DATA <= x"1bfe";
            when "11" & x"fd4" => DATA <= x"fe00";
            when "11" & x"fd5" => DATA <= x"382f";
            when "11" & x"fd6" => DATA <= x"fc01";
            when "11" & x"fd7" => DATA <= x"ffe0";
            when "11" & x"fd8" => DATA <= x"07f8";
            when "11" & x"fd9" => DATA <= x"0c0f";
            when "11" & x"fda" => DATA <= x"41f4";
            when "11" & x"fdb" => DATA <= x"7e00";
            when "11" & x"fdc" => DATA <= x"1fbf";
            when "11" & x"fdd" => DATA <= x"dfcf";
            when "11" & x"fde" => DATA <= x"c783";
            when "11" & x"fdf" => DATA <= x"8189";
            when "11" & x"fe0" => DATA <= x"4017";
            when "11" & x"fe1" => DATA <= x"fe00";
            when "11" & x"fe2" => DATA <= x"785f";
            when "11" & x"fe3" => DATA <= x"f803";
            when "11" & x"fe4" => DATA <= x"ffc0";
            when "11" & x"fe5" => DATA <= x"0ff6";
            when "11" & x"fe6" => DATA <= x"0004";
            when "11" & x"fe7" => DATA <= x"060f";
            when "11" & x"fe8" => DATA <= x"0f8f";
            when "11" & x"fe9" => DATA <= x"c01d";
            when "11" & x"fea" => DATA <= x"fefe";
            when "11" & x"feb" => DATA <= x"7c3c";
            when "11" & x"fec" => DATA <= x"5800";
            when "11" & x"fed" => DATA <= x"07f5";
            when "11" & x"fee" => DATA <= x"ff80";
            when "11" & x"fef" => DATA <= x"3ffc";
            when "11" & x"ff0" => DATA <= x"00ff";
            when "11" & x"ff1" => DATA <= x"1fef";
            when "11" & x"ff2" => DATA <= x"f801";
            when "11" & x"ff3" => DATA <= x"fee0";
            when "11" & x"ff4" => DATA <= x"0000";
            when "11" & x"ff5" => DATA <= x"c1e7";
            when "11" & x"ff6" => DATA <= x"f7f8";
            when "11" & x"ff7" => DATA <= x"03bf";
            when "11" & x"ff8" => DATA <= x"df8e";
            when "11" & x"ff9" => DATA <= x"1460";
            when "11" & x"ffa" => DATA <= x"c401";
            when "11" & x"ffb" => DATA <= x"7fef";
            when "11" & x"ffc" => DATA <= x"c003";
            when "11" & x"ffd" => DATA <= x"dedc";
            when "11" & x"ffe" => DATA <= x"4e07";
            when "11" & x"fff" => DATA <= x"b0ff";
            when others => DATA <= (others => '0');
        end case;
    end process;
end RTL;
