library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tuberom_pdp11 is
    port (
        CLK  : in  std_logic;
        ADDR : in  std_logic_vector(9 downto 0);
        DATA : out std_logic_vector(15 downto 0)
        );
end;

architecture RTL of tuberom_pdp11 is

    signal rom_addr : std_logic_vector(11 downto 0);

begin

    p_addr : process(ADDR)
    begin
        rom_addr             <= (others => '0');
        rom_addr(9 downto 0) <= ADDR;
    end process;

    p_rom : process
    begin
        wait until rising_edge(CLK);
        DATA <= (others => '0');
        case rom_addr is
            when x"000" => DATA <= x"0077";
            when x"001" => DATA <= x"0018";
            when x"002" => DATA <= x"500d";
            when x"003" => DATA <= x"5044";
            when x"004" => DATA <= x"3131";
            when x"005" => DATA <= x"5420";
            when x"006" => DATA <= x"4255";
            when x"007" => DATA <= x"2045";
            when x"008" => DATA <= x"3436";
            when x"009" => DATA <= x"204b";
            when x"00a" => DATA <= x"2e30";
            when x"00b" => DATA <= x"3332";
            when x"00c" => DATA <= x"0d20";
            when x"00d" => DATA <= x"000d";
            when x"00e" => DATA <= x"15c6";
            when x"00f" => DATA <= x"f530";
            when x"010" => DATA <= x"17e6";
            when x"011" => DATA <= x"f5fc";
            when x"012" => DATA <= x"09f7";
            when x"013" => DATA <= x"0540";
            when x"014" => DATA <= x"159f";
            when x"015" => DATA <= x"f5f8";
            when x"016" => DATA <= x"15c1";
            when x"017" => DATA <= x"f804";
            when x"018" => DATA <= x"09f7";
            when x"019" => DATA <= x"007e";
            when x"01a" => DATA <= x"09f7";
            when x"01b" => DATA <= x"045c";
            when x"01c" => DATA <= x"00a1";
            when x"01d" => DATA <= x"09f7";
            when x"01e" => DATA <= x"00ea";
            when x"01f" => DATA <= x"17c6";
            when x"020" => DATA <= x"f5f6";
            when x"021" => DATA <= x"15c1";
            when x"022" => DATA <= x"f85a";
            when x"023" => DATA <= x"09f7";
            when x"024" => DATA <= x"0068";
            when x"025" => DATA <= x"09f7";
            when x"026" => DATA <= x"0254";
            when x"027" => DATA <= x"870c";
            when x"028" => DATA <= x"17c0";
            when x"029" => DATA <= x"f862";
            when x"02a" => DATA <= x"09f7";
            when x"02b" => DATA <= x"0060";
            when x"02c" => DATA <= x"01f4";
            when x"02d" => DATA <= x"4450";
            when x"02e" => DATA <= x"3150";
            when x"02f" => DATA <= x"3e31";
            when x"030" => DATA <= x"002a";
            when x"031" => DATA <= x"f530";
            when x"032" => DATA <= x"20a8";
            when x"033" => DATA <= x"00ff";
            when x"034" => DATA <= x"15c0";
            when x"035" => DATA <= x"007e";
            when x"036" => DATA <= x"09f7";
            when x"037" => DATA <= x"01ae";
            when x"038" => DATA <= x"880f";
            when x"039" => DATA <= x"4511";
            when x"03a" => DATA <= x"6373";
            when x"03b" => DATA <= x"7061";
            when x"03c" => DATA <= x"0065";
            when x"03d" => DATA <= x"17c6";
            when x"03e" => DATA <= x"f5f6";
            when x"03f" => DATA <= x"1001";
            when x"040" => DATA <= x"0a81";
            when x"041" => DATA <= x"09f7";
            when x"042" => DATA <= x"0402";
            when x"043" => DATA <= x"09f7";
            when x"044" => DATA <= x"0028";
            when x"045" => DATA <= x"09f7";
            when x"046" => DATA <= x"03fa";
            when x"047" => DATA <= x"01d7";
            when x"048" => DATA <= x"6000";
            when x"049" => DATA <= x"903f";
            when x"04a" => DATA <= x"fd48";
            when x"04b" => DATA <= x"0087";
            when x"04c" => DATA <= x"e5c1";
            when x"04d" => DATA <= x"0002";
            when x"04e" => DATA <= x"9440";
            when x"04f" => DATA <= x"45c0";
            when x"050" => DATA <= x"ff00";
            when x"051" => DATA <= x"9241";
            when x"052" => DATA <= x"45c1";
            when x"053" => DATA <= x"ff00";
            when x"054" => DATA <= x"00c1";
            when x"055" => DATA <= x"5001";
            when x"056" => DATA <= x"0087";
            when x"057" => DATA <= x"09f7";
            when x"058" => DATA <= x"03d0";
            when x"059" => DATA <= x"9440";
            when x"05a" => DATA <= x"02fc";
            when x"05b" => DATA <= x"0087";
            when x"05c" => DATA <= x"1066";
            when x"05d" => DATA <= x"10a6";
            when x"05e" => DATA <= x"10e6";
            when x"05f" => DATA <= x"1126";
            when x"060" => DATA <= x"1166";
            when x"061" => DATA <= x"1185";
            when x"062" => DATA <= x"2157";
            when x"063" => DATA <= x"f500";
            when x"064" => DATA <= x"8602";
            when x"065" => DATA <= x"15c6";
            when x"066" => DATA <= x"f530";
            when x"067" => DATA <= x"1166";
            when x"068" => DATA <= x"17e6";
            when x"069" => DATA <= x"f5f6";
            when x"06a" => DATA <= x"17e6";
            when x"06b" => DATA <= x"f5fc";
            when x"06c" => DATA <= x"09f7";
            when x"06d" => DATA <= x"0018";
            when x"06e" => DATA <= x"159f";
            when x"06f" => DATA <= x"f5fc";
            when x"070" => DATA <= x"159f";
            when x"071" => DATA <= x"f5f6";
            when x"072" => DATA <= x"1386";
            when x"073" => DATA <= x"1585";
            when x"074" => DATA <= x"1584";
            when x"075" => DATA <= x"1583";
            when x"076" => DATA <= x"1582";
            when x"077" => DATA <= x"1581";
            when x"078" => DATA <= x"0a00";
            when x"079" => DATA <= x"0087";
            when x"07a" => DATA <= x"9401";
            when x"07b" => DATA <= x"a057";
            when x"07c" => DATA <= x"0020";
            when x"07d" => DATA <= x"03fc";
            when x"07e" => DATA <= x"a057";
            when x"07f" => DATA <= x"002a";
            when x"080" => DATA <= x"03f9";
            when x"081" => DATA <= x"0ac0";
            when x"082" => DATA <= x"1001";
            when x"083" => DATA <= x"a417";
            when x"084" => DATA <= x"0021";
            when x"085" => DATA <= x"86fd";
            when x"086" => DATA <= x"0ac0";
            when x"087" => DATA <= x"a417";
            when x"088" => DATA <= x"0020";
            when x"089" => DATA <= x"03fd";
            when x"08a" => DATA <= x"0ac0";
            when x"08b" => DATA <= x"1037";
            when x"08c" => DATA <= x"fcd8";
            when x"08d" => DATA <= x"15c0";
            when x"08e" => DATA <= x"0002";
            when x"08f" => DATA <= x"09f7";
            when x"090" => DATA <= x"051a";
            when x"091" => DATA <= x"09f7";
            when x"092" => DATA <= x"04e6";
            when x"093" => DATA <= x"00b1";
            when x"094" => DATA <= x"09f7";
            when x"095" => DATA <= x"0332";
            when x"096" => DATA <= x"80e2";
            when x"097" => DATA <= x"17c1";
            when x"098" => DATA <= x"f5f8";
            when x"099" => DATA <= x"15c5";
            when x"09a" => DATA <= x"0000";
            when x"09b" => DATA <= x"0c45";
            when x"09c" => DATA <= x"1066";
            when x"09d" => DATA <= x"9c42";
            when x"09e" => DATA <= x"0007";
            when x"09f" => DATA <= x"45c2";
            when x"0a0" => DATA <= x"ff00";
            when x"0a1" => DATA <= x"6081";
            when x"0a2" => DATA <= x"8bd1";
            when x"0a3" => DATA <= x"0226";
            when x"0a4" => DATA <= x"a457";
            when x"0a5" => DATA <= x"0028";
            when x"0a6" => DATA <= x"0223";
            when x"0a7" => DATA <= x"a457";
            when x"0a8" => DATA <= x"0043";
            when x"0a9" => DATA <= x"0220";
            when x"0aa" => DATA <= x"a457";
            when x"0ab" => DATA <= x"0029";
            when x"0ac" => DATA <= x"021d";
            when x"0ad" => DATA <= x"1381";
            when x"0ae" => DATA <= x"9c42";
            when x"0af" => DATA <= x"0006";
            when x"0b0" => DATA <= x"45c2";
            when x"0b1" => DATA <= x"ffb0";
            when x"0b2" => DATA <= x"2097";
            when x"0b3" => DATA <= x"0047";
            when x"0b4" => DATA <= x"0247";
            when x"0b5" => DATA <= x"9c42";
            when x"0b6" => DATA <= x"0006";
            when x"0b7" => DATA <= x"35c2";
            when x"0b8" => DATA <= x"0020";
            when x"0b9" => DATA <= x"030e";
            when x"0ba" => DATA <= x"9c42";
            when x"0bb" => DATA <= x"0007";
            when x"0bc" => DATA <= x"45c2";
            when x"0bd" => DATA <= x"ff00";
            when x"0be" => DATA <= x"6081";
            when x"0bf" => DATA <= x"0a81";
            when x"0c0" => DATA <= x"8bd1";
            when x"0c1" => DATA <= x"02fe";
            when x"0c2" => DATA <= x"65c1";
            when x"0c3" => DATA <= x"0004";
            when x"0c4" => DATA <= x"09f7";
            when x"0c5" => DATA <= x"ff10";
            when x"0c6" => DATA <= x"6581";
            when x"0c7" => DATA <= x"1066";
            when x"0c8" => DATA <= x"55c5";
            when x"0c9" => DATA <= x"0002";
            when x"0ca" => DATA <= x"1581";
            when x"0cb" => DATA <= x"45c1";
            when x"0cc" => DATA <= x"0001";
            when x"0cd" => DATA <= x"1242";
            when x"0ce" => DATA <= x"2097";
            when x"0cf" => DATA <= x"0105";
            when x"0d0" => DATA <= x"871a";
            when x"0d1" => DATA <= x"2097";
            when x"0d2" => DATA <= x"0109";
            when x"0d3" => DATA <= x"8617";
            when x"0d4" => DATA <= x"0bd1";
            when x"0d5" => DATA <= x"1443";
            when x"0d6" => DATA <= x"1444";
            when x"0d7" => DATA <= x"6103";
            when x"0d8" => DATA <= x"1444";
            when x"0d9" => DATA <= x"17c2";
            when x"0da" => DATA <= x"f5f4";
            when x"0db" => DATA <= x"65c1";
            when x"0dc" => DATA <= x"0008";
            when x"0dd" => DATA <= x"0c83";
            when x"0de" => DATA <= x"1452";
            when x"0df" => DATA <= x"0ac3";
            when x"0e0" => DATA <= x"02fd";
            when x"0e1" => DATA <= x"0c84";
            when x"0e2" => DATA <= x"0303";
            when x"0e3" => DATA <= x"0a12";
            when x"0e4" => DATA <= x"0ac4";
            when x"0e5" => DATA <= x"02fd";
            when x"0e6" => DATA <= x"17c1";
            when x"0e7" => DATA <= x"f5f4";
            when x"0e8" => DATA <= x"0a26";
            when x"0e9" => DATA <= x"0a26";
            when x"0ea" => DATA <= x"0a26";
            when x"0eb" => DATA <= x"1066";
            when x"0ec" => DATA <= x"1140";
            when x"0ed" => DATA <= x"15c5";
            when x"0ee" => DATA <= x"0bbc";
            when x"0ef" => DATA <= x"0a04";
            when x"0f0" => DATA <= x"0a03";
            when x"0f1" => DATA <= x"0a02";
            when x"0f2" => DATA <= x"17c1";
            when x"0f3" => DATA <= x"f5f2";
            when x"0f4" => DATA <= x"0c80";
            when x"0f5" => DATA <= x"0305";
            when x"0f6" => DATA <= x"139f";
            when x"0f7" => DATA <= x"f5fc";
            when x"0f8" => DATA <= x"8002";
            when x"0f9" => DATA <= x"139f";
            when x"0fa" => DATA <= x"f5f6";
            when x"0fb" => DATA <= x"0087";
            when x"0fc" => DATA <= x"0c85";
            when x"0fd" => DATA <= x"860b";
            when x"0fe" => DATA <= x"09f7";
            when x"0ff" => DATA <= x"039c";
            when x"100" => DATA <= x"880f";
            when x"101" => DATA <= x"4ef9";
            when x"102" => DATA <= x"746f";
            when x"103" => DATA <= x"5020";
            when x"104" => DATA <= x"5044";
            when x"105" => DATA <= x"3131";
            when x"106" => DATA <= x"6320";
            when x"107" => DATA <= x"646f";
            when x"108" => DATA <= x"0065";
            when x"109" => DATA <= x"0077";
            when x"10a" => DATA <= x"fe28";
            when x"10b" => DATA <= x"15f7";
            when x"10c" => DATA <= x"f804";
            when x"10d" => DATA <= x"fbd6";
            when x"10e" => DATA <= x"0184";
            when x"10f" => DATA <= x"1026";
            when x"110" => DATA <= x"8bc0";
            when x"111" => DATA <= x"810b";
            when x"112" => DATA <= x"15c0";
            when x"113" => DATA <= x"0004";
            when x"114" => DATA <= x"09f7";
            when x"115" => DATA <= x"040a";
            when x"116" => DATA <= x"1380";
            when x"117" => DATA <= x"09f7";
            when x"118" => DATA <= x"040a";
            when x"119" => DATA <= x"09f7";
            when x"11a" => DATA <= x"0228";
            when x"11b" => DATA <= x"1001";
            when x"11c" => DATA <= x"0132";
            when x"11d" => DATA <= x"2017";
            when x"11e" => DATA <= x"0082";
            when x"11f" => DATA <= x"8704";
            when x"120" => DATA <= x"0325";
            when x"121" => DATA <= x"2017";
            when x"122" => DATA <= x"0085";
            when x"123" => DATA <= x"8724";
            when x"124" => DATA <= x"15c0";
            when x"125" => DATA <= x"0006";
            when x"126" => DATA <= x"09f7";
            when x"127" => DATA <= x"03e6";
            when x"128" => DATA <= x"1080";
            when x"129" => DATA <= x"09f7";
            when x"12a" => DATA <= x"03e6";
            when x"12b" => DATA <= x"1580";
            when x"12c" => DATA <= x"09f7";
            when x"12d" => DATA <= x"03e0";
            when x"12e" => DATA <= x"2017";
            when x"12f" => DATA <= x"009d";
            when x"130" => DATA <= x"031f";
            when x"131" => DATA <= x"2017";
            when x"132" => DATA <= x"008e";
            when x"133" => DATA <= x"03d7";
            when x"134" => DATA <= x"1026";
            when x"135" => DATA <= x"09f7";
            when x"136" => DATA <= x"01f0";
            when x"137" => DATA <= x"65c0";
            when x"138" => DATA <= x"ff80";
            when x"139" => DATA <= x"09f7";
            when x"13a" => DATA <= x"01e8";
            when x"13b" => DATA <= x"45c0";
            when x"13c" => DATA <= x"ff00";
            when x"13d" => DATA <= x"1002";
            when x"13e" => DATA <= x"00c0";
            when x"13f" => DATA <= x"1001";
            when x"140" => DATA <= x"09f7";
            when x"141" => DATA <= x"01da";
            when x"142" => DATA <= x"45c0";
            when x"143" => DATA <= x"ff00";
            when x"144" => DATA <= x"5001";
            when x"145" => DATA <= x"0109";
            when x"146" => DATA <= x"15c0";
            when x"147" => DATA <= x"0086";
            when x"148" => DATA <= x"0cc0";
            when x"149" => DATA <= x"1c01";
            when x"14a" => DATA <= x"f4ee";
            when x"14b" => DATA <= x"1042";
            when x"14c" => DATA <= x"00c2";
            when x"14d" => DATA <= x"45c2";
            when x"14e" => DATA <= x"ff00";
            when x"14f" => DATA <= x"1580";
            when x"150" => DATA <= x"0087";
            when x"151" => DATA <= x"0bc0";
            when x"152" => DATA <= x"034d";
            when x"153" => DATA <= x"10e6";
            when x"154" => DATA <= x"10a6";
            when x"155" => DATA <= x"1026";
            when x"156" => DATA <= x"15c0";
            when x"157" => DATA <= x"0008";
            when x"158" => DATA <= x"09f7";
            when x"159" => DATA <= x"0388";
            when x"15a" => DATA <= x"1380";
            when x"15b" => DATA <= x"09f7";
            when x"15c" => DATA <= x"0382";
            when x"15d" => DATA <= x"8bc0";
            when x"15e" => DATA <= x"8003";
            when x"15f" => DATA <= x"9442";
            when x"160" => DATA <= x"9243";
            when x"161" => DATA <= x"010c";
            when x"162" => DATA <= x"15c2";
            when x"163" => DATA <= x"0010";
            when x"164" => DATA <= x"15c3";
            when x"165" => DATA <= x"0010";
            when x"166" => DATA <= x"2017";
            when x"167" => DATA <= x"0015";
            when x"168" => DATA <= x"8605";
            when x"169" => DATA <= x"6000";
            when x"16a" => DATA <= x"65c0";
            when x"16b" => DATA <= x"fb16";
            when x"16c" => DATA <= x"9402";
            when x"16d" => DATA <= x"9203";
            when x"16e" => DATA <= x"1080";
            when x"16f" => DATA <= x"09f7";
            when x"170" => DATA <= x"035a";
            when x"171" => DATA <= x"6081";
            when x"172" => DATA <= x"0ac2";
            when x"173" => DATA <= x"2097";
            when x"174" => DATA <= x"0080";
            when x"175" => DATA <= x"8605";
            when x"176" => DATA <= x"9840";
            when x"177" => DATA <= x"09f7";
            when x"178" => DATA <= x"034a";
            when x"179" => DATA <= x"0ac2";
            when x"17a" => DATA <= x"80fb";
            when x"17b" => DATA <= x"10c0";
            when x"17c" => DATA <= x"09f7";
            when x"17d" => DATA <= x"0340";
            when x"17e" => DATA <= x"60c1";
            when x"17f" => DATA <= x"0ac3";
            when x"180" => DATA <= x"20d7";
            when x"181" => DATA <= x"0080";
            when x"182" => DATA <= x"8605";
            when x"183" => DATA <= x"09f7";
            when x"184" => DATA <= x"0154";
            when x"185" => DATA <= x"9021";
            when x"186" => DATA <= x"0ac3";
            when x"187" => DATA <= x"80fb";
            when x"188" => DATA <= x"1580";
            when x"189" => DATA <= x"1582";
            when x"18a" => DATA <= x"1583";
            when x"18b" => DATA <= x"0087";
            when x"18c" => DATA <= x"0500";
            when x"18d" => DATA <= x"0005";
            when x"18e" => DATA <= x"0500";
            when x"18f" => DATA <= x"0005";
            when x"190" => DATA <= x"0504";
            when x"191" => DATA <= x"0005";
            when x"192" => DATA <= x"0008";
            when x"193" => DATA <= x"000e";
            when x"194" => DATA <= x"0504";
            when x"195" => DATA <= x"0901";
            when x"196" => DATA <= x"0501";
            when x"197" => DATA <= x"0005";
            when x"198" => DATA <= x"0800";
            when x"199" => DATA <= x"1910";
            when x"19a" => DATA <= x"0020";
            when x"19b" => DATA <= x"0110";
            when x"19c" => DATA <= x"0d0d";
            when x"19d" => DATA <= x"8000";
            when x"19e" => DATA <= x"0808";
            when x"19f" => DATA <= x"8080";
            when x"1a0" => DATA <= x"15c0";
            when x"1a1" => DATA <= x"000a";
            when x"1a2" => DATA <= x"09f7";
            when x"1a3" => DATA <= x"02f4";
            when x"1a4" => DATA <= x"65c1";
            when x"1a5" => DATA <= x"0002";
            when x"1a6" => DATA <= x"15c2";
            when x"1a7" => DATA <= x"0003";
            when x"1a8" => DATA <= x"09f7";
            when x"1a9" => DATA <= x"02c6";
            when x"1aa" => DATA <= x"15c0";
            when x"1ab" => DATA <= x"0007";
            when x"1ac" => DATA <= x"09f7";
            when x"1ad" => DATA <= x"02e0";
            when x"1ae" => DATA <= x"0a00";
            when x"1af" => DATA <= x"09f7";
            when x"1b0" => DATA <= x"02da";
            when x"1b1" => DATA <= x"09f7";
            when x"1b2" => DATA <= x"00f8";
            when x"1b3" => DATA <= x"65c0";
            when x"1b4" => DATA <= x"ff80";
            when x"1b5" => DATA <= x"870b";
            when x"1b6" => DATA <= x"09f7";
            when x"1b7" => DATA <= x"fd28";
            when x"1b8" => DATA <= x"0a02";
            when x"1b9" => DATA <= x"09f7";
            when x"1ba" => DATA <= x"00e8";
            when x"1bb" => DATA <= x"9011";
            when x"1bc" => DATA <= x"0a82";
            when x"1bd" => DATA <= x"2017";
            when x"1be" => DATA <= x"000d";
            when x"1bf" => DATA <= x"02f9";
            when x"1c0" => DATA <= x"0ac2";
            when x"1c1" => DATA <= x"0087";
            when x"1c2" => DATA <= x"10a6";
            when x"1c3" => DATA <= x"1066";
            when x"1c4" => DATA <= x"1026";
            when x"1c5" => DATA <= x"15c0";
            when x"1c6" => DATA <= x"000c";
            when x"1c7" => DATA <= x"09f7";
            when x"1c8" => DATA <= x"02a4";
            when x"1c9" => DATA <= x"1081";
            when x"1ca" => DATA <= x"15c2";
            when x"1cb" => DATA <= x"0004";
            when x"1cc" => DATA <= x"09f7";
            when x"1cd" => DATA <= x"027e";
            when x"1ce" => DATA <= x"1580";
            when x"1cf" => DATA <= x"09f7";
            when x"1d0" => DATA <= x"029a";
            when x"1d1" => DATA <= x"09f7";
            when x"1d2" => DATA <= x"00b8";
            when x"1d3" => DATA <= x"1026";
            when x"1d4" => DATA <= x"15c2";
            when x"1d5" => DATA <= x"0004";
            when x"1d6" => DATA <= x"0133";
            when x"1d7" => DATA <= x"1026";
            when x"1d8" => DATA <= x"15c0";
            when x"1d9" => DATA <= x"0012";
            when x"1da" => DATA <= x"09f7";
            when x"1db" => DATA <= x"0284";
            when x"1dc" => DATA <= x"1580";
            when x"1dd" => DATA <= x"09f7";
            when x"1de" => DATA <= x"027e";
            when x"1df" => DATA <= x"0bc0";
            when x"1e0" => DATA <= x"0206";
            when x"1e1" => DATA <= x"09f7";
            when x"1e2" => DATA <= x"0274";
            when x"1e3" => DATA <= x"09f7";
            when x"1e4" => DATA <= x"0094";
            when x"1e5" => DATA <= x"0a00";
            when x"1e6" => DATA <= x"0087";
            when x"1e7" => DATA <= x"1066";
            when x"1e8" => DATA <= x"09f7";
            when x"1e9" => DATA <= x"0238";
            when x"1ea" => DATA <= x"09f7";
            when x"1eb" => DATA <= x"0086";
            when x"1ec" => DATA <= x"1581";
            when x"1ed" => DATA <= x"0087";
            when x"1ee" => DATA <= x"10a6";
            when x"1ef" => DATA <= x"1066";
            when x"1f0" => DATA <= x"1026";
            when x"1f1" => DATA <= x"15c0";
            when x"1f2" => DATA <= x"0014";
            when x"1f3" => DATA <= x"09f7";
            when x"1f4" => DATA <= x"0252";
            when x"1f5" => DATA <= x"65c1";
            when x"1f6" => DATA <= x"0002";
            when x"1f7" => DATA <= x"15c2";
            when x"1f8" => DATA <= x"0010";
            when x"1f9" => DATA <= x"09f7";
            when x"1fa" => DATA <= x"0224";
            when x"1fb" => DATA <= x"09f7";
            when x"1fc" => DATA <= x"fc9e";
            when x"1fd" => DATA <= x"09f7";
            when x"1fe" => DATA <= x"020e";
            when x"1ff" => DATA <= x"1580";
            when x"200" => DATA <= x"09f7";
            when x"201" => DATA <= x"0238";
            when x"202" => DATA <= x"09f7";
            when x"203" => DATA <= x"0056";
            when x"204" => DATA <= x"1381";
            when x"205" => DATA <= x"1026";
            when x"206" => DATA <= x"65c1";
            when x"207" => DATA <= x"0002";
            when x"208" => DATA <= x"15c2";
            when x"209" => DATA <= x"0010";
            when x"20a" => DATA <= x"09f7";
            when x"20b" => DATA <= x"0210";
            when x"20c" => DATA <= x"1580";
            when x"20d" => DATA <= x"1581";
            when x"20e" => DATA <= x"1582";
            when x"20f" => DATA <= x"0087";
            when x"210" => DATA <= x"10a6";
            when x"211" => DATA <= x"1026";
            when x"212" => DATA <= x"15c0";
            when x"213" => DATA <= x"0016";
            when x"214" => DATA <= x"09f7";
            when x"215" => DATA <= x"0210";
            when x"216" => DATA <= x"15c2";
            when x"217" => DATA <= x"000d";
            when x"218" => DATA <= x"09f7";
            when x"219" => DATA <= x"01e6";
            when x"21a" => DATA <= x"1580";
            when x"21b" => DATA <= x"09f7";
            when x"21c" => DATA <= x"0202";
            when x"21d" => DATA <= x"15c2";
            when x"21e" => DATA <= x"000d";
            when x"21f" => DATA <= x"09f7";
            when x"220" => DATA <= x"01e6";
            when x"221" => DATA <= x"1582";
            when x"222" => DATA <= x"0108";
            when x"223" => DATA <= x"15c0";
            when x"224" => DATA <= x"000e";
            when x"225" => DATA <= x"09f7";
            when x"226" => DATA <= x"01e8";
            when x"227" => DATA <= x"0103";
            when x"228" => DATA <= x"0a00";
            when x"229" => DATA <= x"09f7";
            when x"22a" => DATA <= x"01e6";
            when x"22b" => DATA <= x"09f7";
            when x"22c" => DATA <= x"0004";
            when x"22d" => DATA <= x"65c0";
            when x"22e" => DATA <= x"ff80";
            when x"22f" => DATA <= x"97c0";
            when x"230" => DATA <= x"fff4";
            when x"231" => DATA <= x"80fd";
            when x"232" => DATA <= x"97c0";
            when x"233" => DATA <= x"fff6";
            when x"234" => DATA <= x"0087";
            when x"235" => DATA <= x"1026";
            when x"236" => DATA <= x"15c0";
            when x"237" => DATA <= x"0010";
            when x"238" => DATA <= x"09f7";
            when x"239" => DATA <= x"01c2";
            when x"23a" => DATA <= x"1380";
            when x"23b" => DATA <= x"09f7";
            when x"23c" => DATA <= x"01c2";
            when x"23d" => DATA <= x"09f7";
            when x"23e" => DATA <= x"ffe0";
            when x"23f" => DATA <= x"1580";
            when x"240" => DATA <= x"0087";
            when x"241" => DATA <= x"25c0";
            when x"242" => DATA <= x"000d";
            when x"243" => DATA <= x"0206";
            when x"244" => DATA <= x"15c0";
            when x"245" => DATA <= x"000a";
            when x"246" => DATA <= x"09f7";
            when x"247" => DATA <= x"0004";
            when x"248" => DATA <= x"15c0";
            when x"249" => DATA <= x"000d";
            when x"24a" => DATA <= x"35df";
            when x"24b" => DATA <= x"0040";
            when x"24c" => DATA <= x"fff0";
            when x"24d" => DATA <= x"03fc";
            when x"24e" => DATA <= x"901f";
            when x"24f" => DATA <= x"fff2";
            when x"250" => DATA <= x"0087";
            when x"251" => DATA <= x"880f";
            when x"252" => DATA <= x"42ff";
            when x"253" => DATA <= x"6461";
            when x"254" => DATA <= x"0000";
            when x"255" => DATA <= x"45f6";
            when x"256" => DATA <= x"fff0";
            when x"257" => DATA <= x"0002";
            when x"258" => DATA <= x"17e6";
            when x"259" => DATA <= x"f5e0";
            when x"25a" => DATA <= x"17e6";
            when x"25b" => DATA <= x"f5ec";
            when x"25c" => DATA <= x"119f";
            when x"25d" => DATA <= x"f5ec";
            when x"25e" => DATA <= x"15df";
            when x"25f" => DATA <= x"fce0";
            when x"260" => DATA <= x"f5e0";
            when x"261" => DATA <= x"0be6";
            when x"262" => DATA <= x"1026";
            when x"263" => DATA <= x"1d80";
            when x"264" => DATA <= x"0008";
            when x"265" => DATA <= x"1800";
            when x"266" => DATA <= x"45c0";
            when x"267" => DATA <= x"ff00";
            when x"268" => DATA <= x"6000";
            when x"269" => DATA <= x"67c0";
            when x"26a" => DATA <= x"f5ee";
            when x"26b" => DATA <= x"1236";
            when x"26c" => DATA <= x"0002";
            when x"26d" => DATA <= x"1580";
            when x"26e" => DATA <= x"09de";
            when x"26f" => DATA <= x"8405";
            when x"270" => DATA <= x"17c6";
            when x"271" => DATA <= x"f5ec";
            when x"272" => DATA <= x"55f6";
            when x"273" => DATA <= x"0002";
            when x"274" => DATA <= x"0006";
            when x"275" => DATA <= x"8603";
            when x"276" => DATA <= x"55f6";
            when x"277" => DATA <= x"0001";
            when x"278" => DATA <= x"0006";
            when x"279" => DATA <= x"159f";
            when x"27a" => DATA <= x"f5ec";
            when x"27b" => DATA <= x"159f";
            when x"27c" => DATA <= x"f5e0";
            when x"27d" => DATA <= x"0002";
            when x"27e" => DATA <= x"1d80";
            when x"27f" => DATA <= x"0006";
            when x"280" => DATA <= x"1db6";
            when x"281" => DATA <= x"0004";
            when x"282" => DATA <= x"0006";
            when x"283" => DATA <= x"0087";
            when x"284" => DATA <= x"0bd6";
            when x"285" => DATA <= x"159f";
            when x"286" => DATA <= x"f5ec";
            when x"287" => DATA <= x"159f";
            when x"288" => DATA <= x"f5e0";
            when x"289" => DATA <= x"1026";
            when x"28a" => DATA <= x"810b";
            when x"28b" => DATA <= x"2017";
            when x"28c" => DATA <= x"0100";
            when x"28d" => DATA <= x"861b";
            when x"28e" => DATA <= x"6000";
            when x"28f" => DATA <= x"67c0";
            when x"290" => DATA <= x"f5ee";
            when x"291" => DATA <= x"1226";
            when x"292" => DATA <= x"0bc1";
            when x"293" => DATA <= x"0314";
            when x"294" => DATA <= x"1048";
            when x"295" => DATA <= x"0112";
            when x"296" => DATA <= x"0a40";
            when x"297" => DATA <= x"2017";
            when x"298" => DATA <= x"000a";
            when x"299" => DATA <= x"860f";
            when x"29a" => DATA <= x"6000";
            when x"29b" => DATA <= x"6000";
            when x"29c" => DATA <= x"65c0";
            when x"29d" => DATA <= x"f5d8";
            when x"29e" => DATA <= x"1226";
            when x"29f" => DATA <= x"0bc1";
            when x"2a0" => DATA <= x"0301"; -- was 17f6
            when x"2a1" => DATA <= x"1048"; -- was f5e0
            when x"2a2" => DATA <= x"0bd0";
            when x"2a3" => DATA <= x"1226";
            when x"2a4" => DATA <= x"0bc2";
            when x"2a5" => DATA <= x"0301";
            when x"2a6" => DATA <= x"1088";
            when x"2a7" => DATA <= x"1582";
            when x"2a8" => DATA <= x"1581";
            when x"2a9" => DATA <= x"1580";
            when x"2aa" => DATA <= x"0002";
            when x"2ab" => DATA <= x"0bc0";
            when x"2ac" => DATA <= x"0304";
            when x"2ad" => DATA <= x"2017";
            when x"2ae" => DATA <= x"0003";
            when x"2af" => DATA <= x"871d";
            when x"2b0" => DATA <= x"0303";
            when x"2b1" => DATA <= x"0087";
            when x"2b2" => DATA <= x"007f";
            when x"2b3" => DATA <= x"f870";
            when x"2b4" => DATA <= x"0a00";
            when x"2b5" => DATA <= x"15d0";
            when x"2b6" => DATA <= x"ff92";
            when x"2b7" => DATA <= x"0a10";
            when x"2b8" => DATA <= x"2017";
            when x"2b9" => DATA <= x"0100";
            when x"2ba" => DATA <= x"02fa";
            when x"2bb" => DATA <= x"15df";
            when x"2bc" => DATA <= x"fca2";
            when x"2bd" => DATA <= x"001c";
            when x"2be" => DATA <= x"15df";
            when x"2bf" => DATA <= x"fcaa";
            when x"2c0" => DATA <= x"0018";
            when x"2c1" => DATA <= x"15df";
            when x"2c2" => DATA <= x"ff8e";
            when x"2c3" => DATA <= x"0080";
            when x"2c4" => DATA <= x"15df";
            when x"2c5" => DATA <= x"00e0";
            when x"2c6" => DATA <= x"0082";
            when x"2c7" => DATA <= x"15df";
            when x"2c8" => DATA <= x"fe62";
            when x"2c9" => DATA <= x"0084";
            when x"2ca" => DATA <= x"15df";
            when x"2cb" => DATA <= x"00c0";
            when x"2cc" => DATA <= x"0086";
            when x"2cd" => DATA <= x"0c00";
            when x"2ce" => DATA <= x"15c0";
            when x"2cf" => DATA <= x"000c";
            when x"2d0" => DATA <= x"15c1";
            when x"2d1" => DATA <= x"fdc2";
            when x"2d2" => DATA <= x"15c2";
            when x"2d3" => DATA <= x"f5d8";
            when x"2d4" => DATA <= x"8702";
            when x"2d5" => DATA <= x"65c0";
            when x"2d6" => DATA <= x"0018";
            when x"2d7" => DATA <= x"1452";
            when x"2d8" => DATA <= x"0ac0";
            when x"2d9" => DATA <= x"02fd";
            when x"2da" => DATA <= x"8705";
            when x"2db" => DATA <= x"15c0";
            when x"2dc" => DATA <= x"00f0";
            when x"2dd" => DATA <= x"1252";
            when x"2de" => DATA <= x"0ac0";
            when x"2df" => DATA <= x"02fd";
            when x"2e0" => DATA <= x"0087";
            when x"2e1" => DATA <= x"f83e";
            when x"2e2" => DATA <= x"0000";
            when x"2e3" => DATA <= x"f890";
            when x"2e4" => DATA <= x"f5ff";
            when x"2e5" => DATA <= x"f87a";
            when x"2e6" => DATA <= x"f500";
            when x"2e7" => DATA <= x"fd62";
            when x"2e8" => DATA <= x"0000";
            when x"2e9" => DATA <= x"ff92";
            when x"2ea" => DATA <= x"0000";
            when x"2eb" => DATA <= x"0000";
            when x"2ec" => DATA <= x"f600";
            when x"2ed" => DATA <= x"0000";
            when x"2ee" => DATA <= x"f804";
            when x"2ef" => DATA <= x"0100";
            when x"2f0" => DATA <= x"f500";
            when x"2f1" => DATA <= x"f83e";
            when x"2f2" => DATA <= x"0000";
            when x"2f3" => DATA <= x"f83e";
            when x"2f4" => DATA <= x"0000";
            when x"2f5" => DATA <= x"fd64";
            when x"2f6" => DATA <= x"f8b8";
            when x"2f7" => DATA <= x"fa1e";
            when x"2f8" => DATA <= x"faa2";
            when x"2f9" => DATA <= x"fc94";
            when x"2fa" => DATA <= x"fc88";
            when x"2fb" => DATA <= x"fc50";
            when x"2fc" => DATA <= x"fbdc";
            when x"2fd" => DATA <= x"fb84";
            when x"2fe" => DATA <= x"fc46";
            when x"2ff" => DATA <= x"fc6a";
            when x"300" => DATA <= x"fc20";
            when x"301" => DATA <= x"fbae";
            when x"302" => DATA <= x"fd56";
            when x"303" => DATA <= x"fd08";
            when x"304" => DATA <= x"fcfc";
            when x"305" => DATA <= x"fd62";
            when x"306" => DATA <= x"9440";
            when x"307" => DATA <= x"09f7";
            when x"308" => DATA <= x"002a";
            when x"309" => DATA <= x"2017";
            when x"30a" => DATA <= x"000d";
            when x"30b" => DATA <= x"02fa";
            when x"30c" => DATA <= x"0087";
            when x"30d" => DATA <= x"6081";
            when x"30e" => DATA <= x"9840";
            when x"30f" => DATA <= x"09f7";
            when x"310" => DATA <= x"001a";
            when x"311" => DATA <= x"0ac2";
            when x"312" => DATA <= x"02fb";
            when x"313" => DATA <= x"0087";
            when x"314" => DATA <= x"6081";
            when x"315" => DATA <= x"09f7";
            when x"316" => DATA <= x"fe30";
            when x"317" => DATA <= x"9021";
            when x"318" => DATA <= x"0ac2";
            when x"319" => DATA <= x"02fb";
            when x"31a" => DATA <= x"0087";
            when x"31b" => DATA <= x"09f7";
            when x"31c" => DATA <= x"0002";
            when x"31d" => DATA <= x"1040";
            when x"31e" => DATA <= x"35df";
            when x"31f" => DATA <= x"0040";
            when x"320" => DATA <= x"fff4";
            when x"321" => DATA <= x"03fc";
            when x"322" => DATA <= x"901f";
            when x"323" => DATA <= x"fff6";
            when x"324" => DATA <= x"0087";
            when x"325" => DATA <= x"97c0";
            when x"326" => DATA <= x"fff0";
            when x"327" => DATA <= x"80fd";
            when x"328" => DATA <= x"97c0";
            when x"329" => DATA <= x"fff2";
            when x"32a" => DATA <= x"0087";
            when x"32b" => DATA <= x"97c0";
            when x"32c" => DATA <= x"fffc";
            when x"32d" => DATA <= x"80fd";
            when x"32e" => DATA <= x"97c0";
            when x"32f" => DATA <= x"fffe";
            when x"330" => DATA <= x"0087";
            when x"331" => DATA <= x"1026";
            when x"332" => DATA <= x"97c0";
            when x"333" => DATA <= x"fffc";
            when x"334" => DATA <= x"811c";
            when x"335" => DATA <= x"97c0";
            when x"336" => DATA <= x"fff0";
            when x"337" => DATA <= x"8103";
            when x"338" => DATA <= x"1580";
            when x"339" => DATA <= x"007f";
            when x"33a" => DATA <= x"f772";
            when x"33b" => DATA <= x"97c0";
            when x"33c" => DATA <= x"fff2";
            when x"33d" => DATA <= x"8110";
            when x"33e" => DATA <= x"1066";
            when x"33f" => DATA <= x"10a6";
            when x"340" => DATA <= x"09f7";
            when x"341" => DATA <= x"ffc6";
            when x"342" => DATA <= x"1002";
            when x"343" => DATA <= x"09f7";
            when x"344" => DATA <= x"ffc0";
            when x"345" => DATA <= x"1001";
            when x"346" => DATA <= x"09f7";
            when x"347" => DATA <= x"ffba";
            when x"348" => DATA <= x"09ff";
            when x"349" => DATA <= x"f750";
            when x"34a" => DATA <= x"1582";
            when x"34b" => DATA <= x"1581";
            when x"34c" => DATA <= x"1580";
            when x"34d" => DATA <= x"0002";
            when x"34e" => DATA <= x"09ff";
            when x"34f" => DATA <= x"f73c";
            when x"350" => DATA <= x"0156";
            when x"351" => DATA <= x"97c0";
            when x"352" => DATA <= x"fffe";
            when x"353" => DATA <= x"8013";
            when x"354" => DATA <= x"1066";
            when x"355" => DATA <= x"09f7";
            when x"356" => DATA <= x"fdb0";
            when x"357" => DATA <= x"17c1";
            when x"358" => DATA <= x"f5e2";
            when x"359" => DATA <= x"09f7";
            when x"35a" => DATA <= x"fda8";
            when x"35b" => DATA <= x"9011";
            when x"35c" => DATA <= x"09f7";
            when x"35d" => DATA <= x"fda2";
            when x"35e" => DATA <= x"9011";
            when x"35f" => DATA <= x"02fc";
            when x"360" => DATA <= x"1581";
            when x"361" => DATA <= x"1580";
            when x"362" => DATA <= x"17c0";
            when x"363" => DATA <= x"f5e2";
            when x"364" => DATA <= x"17ce";
            when x"365" => DATA <= x"f5e0";
            when x"366" => DATA <= x"0002";
            when x"367" => DATA <= x"1066";
            when x"368" => DATA <= x"1001";
            when x"369" => DATA <= x"09f7";
            when x"36a" => DATA <= x"ff80";
            when x"36b" => DATA <= x"2057";
            when x"36c" => DATA <= x"0005";
            when x"36d" => DATA <= x"03dd";
            when x"36e" => DATA <= x"09f7";
            when x"36f" => DATA <= x"ff76";
            when x"370" => DATA <= x"901f";
            when x"371" => DATA <= x"f5fb";
            when x"372" => DATA <= x"09f7";
            when x"373" => DATA <= x"ff6e";
            when x"374" => DATA <= x"901f";
            when x"375" => DATA <= x"f5fa";
            when x"376" => DATA <= x"09f7";
            when x"377" => DATA <= x"ff66";
            when x"378" => DATA <= x"901f";
            when x"379" => DATA <= x"f5f9";
            when x"37a" => DATA <= x"09f7";
            when x"37b" => DATA <= x"ff5e";
            when x"37c" => DATA <= x"901f";
            when x"37d" => DATA <= x"f5f8";
            when x"37e" => DATA <= x"97c0";
            when x"37f" => DATA <= x"fffa";
            when x"380" => DATA <= x"97c0";
            when x"381" => DATA <= x"fffa";
            when x"382" => DATA <= x"09f7";
            when x"383" => DATA <= x"ff4e";
            when x"384" => DATA <= x"6041";
            when x"385" => DATA <= x"1c5f";
            when x"386" => DATA <= x"ff94";
            when x"387" => DATA <= x"0080";
            when x"388" => DATA <= x"17c0";
            when x"389" => DATA <= x"f5f8";
            when x"38a" => DATA <= x"2057";
            when x"38b" => DATA <= x"000c";
            when x"38c" => DATA <= x"87be";
            when x"38d" => DATA <= x"030a";
            when x"38e" => DATA <= x"15c1";
            when x"38f" => DATA <= x"0100";
            when x"390" => DATA <= x"8bdf";
            when x"391" => DATA <= x"fff8";
            when x"392" => DATA <= x"80fd";
            when x"393" => DATA <= x"97d0";
            when x"394" => DATA <= x"fffa";
            when x"395" => DATA <= x"0ac1";
            when x"396" => DATA <= x"02f9";
            when x"397" => DATA <= x"010e";
            when x"398" => DATA <= x"15c1";
            when x"399" => DATA <= x"0100";
            when x"39a" => DATA <= x"8bdf";
            when x"39b" => DATA <= x"fff8";
            when x"39c" => DATA <= x"80fd";
            when x"39d" => DATA <= x"941f";
            when x"39e" => DATA <= x"fffa";
            when x"39f" => DATA <= x"0ac1";
            when x"3a0" => DATA <= x"02f9";
            when x"3a1" => DATA <= x"8bdf";
            when x"3a2" => DATA <= x"fff8";
            when x"3a3" => DATA <= x"80fd";
            when x"3a4" => DATA <= x"8a1f";
            when x"3a5" => DATA <= x"fffa";
            when x"3a6" => DATA <= x"1581";
            when x"3a7" => DATA <= x"101f";
            when x"3a8" => DATA <= x"f5f8";
            when x"3a9" => DATA <= x"1580";
            when x"3aa" => DATA <= x"0002";
            when x"3ab" => DATA <= x"1026";
            when x"3ac" => DATA <= x"17c0";
            when x"3ad" => DATA <= x"f5f8";
            when x"3ae" => DATA <= x"97d0";
            when x"3af" => DATA <= x"fffa";
            when x"3b0" => DATA <= x"97d0";
            when x"3b1" => DATA <= x"fffa";
            when x"3b2" => DATA <= x"01f4";
            when x"3b3" => DATA <= x"1026";
            when x"3b4" => DATA <= x"17c0";
            when x"3b5" => DATA <= x"f5f8";
            when x"3b6" => DATA <= x"941f";
            when x"3b7" => DATA <= x"fffa";
            when x"3b8" => DATA <= x"941f";
            when x"3b9" => DATA <= x"fffa";
            when x"3ba" => DATA <= x"01ec";
            when x"3bb" => DATA <= x"1026";
            when x"3bc" => DATA <= x"17c0";
            when x"3bd" => DATA <= x"f5f8";
            when x"3be" => DATA <= x"97d0";
            when x"3bf" => DATA <= x"fffa";
            when x"3c0" => DATA <= x"01e6";
            when x"3c1" => DATA <= x"1026";
            when x"3c2" => DATA <= x"17c0";
            when x"3c3" => DATA <= x"f5f8";
            when x"3c4" => DATA <= x"941f";
            when x"3c5" => DATA <= x"fffa";
            when x"3c6" => DATA <= x"01e0";
            when x"3c7" => DATA <= x"8a1f";
            when x"3c8" => DATA <= x"fffa";
            when x"3c9" => DATA <= x"0002";
            when x"3ca" => DATA <= x"ff82";
            when x"3cb" => DATA <= x"ff76";
            when x"3cc" => DATA <= x"ff66";
            when x"3cd" => DATA <= x"ff56";
            when x"3ce" => DATA <= x"ff8e";
            when x"3cf" => DATA <= x"ff8e";
            when x"3d0" => DATA <= x"ff8e";
            when x"3d1" => DATA <= x"ff8e";
            when x"3d2" => DATA <= x"0000";
            when x"3d3" => DATA <= x"0000";
            when x"3d4" => DATA <= x"0000";
            when x"3d5" => DATA <= x"0000";
            when x"3d6" => DATA <= x"0000";
            when x"3d7" => DATA <= x"0000";
            when x"3d8" => DATA <= x"0000";
            when x"3d9" => DATA <= x"0000";
            when x"3da" => DATA <= x"0000";
            when x"3db" => DATA <= x"0000";
            when x"3dc" => DATA <= x"0000";
            when x"3dd" => DATA <= x"0000";
            when x"3de" => DATA <= x"0000";
            when x"3df" => DATA <= x"0000";
            when x"3e0" => DATA <= x"0000";
            when x"3e1" => DATA <= x"0000";
            when x"3e2" => DATA <= x"0000";
            when x"3e3" => DATA <= x"0000";
            when x"3e4" => DATA <= x"0000";
            when x"3e5" => DATA <= x"0000";
            when x"3e6" => DATA <= x"0000";
            when x"3e7" => DATA <= x"0000";
            when x"3e8" => DATA <= x"0000";
            when x"3e9" => DATA <= x"0000";
            when x"3ea" => DATA <= x"0000";
            when x"3eb" => DATA <= x"0000";
            when x"3ec" => DATA <= x"0000";
            when x"3ed" => DATA <= x"0000";
            when x"3ee" => DATA <= x"0000";
            when x"3ef" => DATA <= x"0000";
            when x"3f0" => DATA <= x"0000";
            when x"3f1" => DATA <= x"0000";
            when x"3f2" => DATA <= x"0000";
            when x"3f3" => DATA <= x"0000";
            when x"3f4" => DATA <= x"0000";
            when x"3f5" => DATA <= x"0000";
            when x"3f6" => DATA <= x"0000";
            when x"3f7" => DATA <= x"0000";
            when x"3f8" => DATA <= x"0000";
            when x"3f9" => DATA <= x"0000";
            when x"3fa" => DATA <= x"0000";
            when x"3fb" => DATA <= x"0000";
            when x"3fc" => DATA <= x"0000";
            when x"3fd" => DATA <= x"0000";
            when x"3fe" => DATA <= x"0000";
            when x"3ff" => DATA <= x"0000";
            when others => DATA <= (others => '0');
        end case;
    end process;
end RTL;
