library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity tuberom_65c102_banner is
    port (
        CLK  : in  std_logic;
        ADDR : in  std_logic_vector(10 downto 0);
        DATA : out std_logic_vector(7 downto 0)
        );
end;

architecture RTL of tuberom_65c102_banner is

    type   ram_type is array (0 to 2047) of std_logic_vector (7 downto 0);

    signal RAM                 : ram_type := (
        16#000# => x"a2",
        16#001# => x"00",
        16#002# => x"bd",
        16#003# => x"00",
        16#004# => x"ff",
        16#005# => x"9d",
        16#006# => x"00",
        16#007# => x"ff",
        16#008# => x"ca",
        16#009# => x"d0",
        16#00a# => x"f7",
        16#00b# => x"a2",
        16#00c# => x"36",
        16#00d# => x"bd",
        16#00e# => x"80",
        16#00f# => x"ff",
        16#010# => x"9d",
        16#011# => x"00",
        16#012# => x"02",
        16#013# => x"ca",
        16#014# => x"10",
        16#015# => x"f7",
        16#016# => x"9a",
        16#017# => x"a2",
        16#018# => x"f0",
        16#019# => x"bd",
        16#01a# => x"ff",
        16#01b# => x"fd",
        16#01c# => x"9d",
        16#01d# => x"ff",
        16#01e# => x"fd",
        16#01f# => x"ca",
        16#020# => x"d0",
        16#021# => x"f7",
        16#022# => x"a0",
        16#023# => x"00",
        16#024# => x"84",
        16#025# => x"f8",
        16#026# => x"a9",
        16#027# => x"f8",
        16#028# => x"85",
        16#029# => x"f9",
        16#02a# => x"b1",
        16#02b# => x"f8",
        16#02c# => x"91",
        16#02d# => x"f8",
        16#02e# => x"c8",
        16#02f# => x"d0",
        16#030# => x"f9",
        16#031# => x"e6",
        16#032# => x"f9",
        16#033# => x"a5",
        16#034# => x"f9",
        16#035# => x"c9",
        16#036# => x"fe",
        16#037# => x"d0",
        16#038# => x"f1",
        16#039# => x"a2",
        16#03a# => x"10",
        16#03b# => x"bd",
        16#03c# => x"59",
        16#03d# => x"f8",
        16#03e# => x"9d",
        16#03f# => x"00",
        16#040# => x"01",
        16#041# => x"ca",
        16#042# => x"10",
        16#043# => x"f7",
        16#044# => x"a5",
        16#045# => x"ee",
        16#046# => x"85",
        16#047# => x"f6",
        16#048# => x"a5",
        16#049# => x"ef",
        16#04a# => x"85",
        16#04b# => x"f7",
        16#04c# => x"a9",
        16#04d# => x"00",
        16#04e# => x"85",
        16#04f# => x"ff",
        16#050# => x"85",
        16#051# => x"f2",
        16#052# => x"a9",
        16#053# => x"f8",
        16#054# => x"85",
        16#055# => x"f3",
        16#056# => x"4c",
        16#057# => x"00",
        16#058# => x"01",
        16#059# => x"ad",
        16#05a# => x"f8",
        16#05b# => x"fe",
        16#05c# => x"58",
        16#05d# => x"4c",
        16#05e# => x"60",
        16#05f# => x"f8",
        16#060# => x"20",
        16#061# => x"a5",
        16#062# => x"fe",
        16#063# => x"0a",
        16#064# => x"41",
        16#065# => x"63",
        16#066# => x"6f",
        16#067# => x"72",
        16#068# => x"6e",
        16#069# => x"20",
        16#06a# => x"54",
        16#06b# => x"55",
        16#06c# => x"42",
        16#06d# => x"45",
        16#06e# => x"20",
        16#06f# => x"3f",
        16#070# => x"3f",
        16#071# => x"4d",
        16#072# => x"48",
        16#073# => x"7a",
        16#074# => x"20",
        16#075# => x"36",
        16#076# => x"35",
        16#077# => x"43",
        16#078# => x"31",
        16#079# => x"30",
        16#07a# => x"32",
        16#07b# => x"20",
        16#07c# => x"43",
        16#07d# => x"6f",
        16#07e# => x"2d",
        16#07f# => x"50",
        16#080# => x"72",
        16#081# => x"6f",
        16#082# => x"0a",
        16#083# => x"0a",
        16#084# => x"0d",
        16#085# => x"00",
        16#086# => x"ea",
        16#087# => x"a9",
        16#088# => x"98",
        16#089# => x"8d",
        16#08a# => x"5e",
        16#08b# => x"f8",
        16#08c# => x"a9",
        16#08d# => x"f8",
        16#08e# => x"8d",
        16#08f# => x"5f",
        16#090# => x"f8",
        16#091# => x"20",
        16#092# => x"80",
        16#093# => x"f9",
        16#094# => x"c9",
        16#095# => x"80",
        16#096# => x"f0",
        16#097# => x"28",
        16#098# => x"a9",
        16#099# => x"2a",
        16#09a# => x"20",
        16#09b# => x"ee",
        16#09c# => x"ff",
        16#09d# => x"a2",
        16#09e# => x"68",
        16#09f# => x"a0",
        16#0a0# => x"f9",
        16#0a1# => x"a9",
        16#0a2# => x"00",
        16#0a3# => x"20",
        16#0a4# => x"f1",
        16#0a5# => x"ff",
        16#0a6# => x"b0",
        16#0a7# => x"0a",
        16#0a8# => x"a2",
        16#0a9# => x"36",
        16#0aa# => x"a0",
        16#0ab# => x"02",
        16#0ac# => x"20",
        16#0ad# => x"f7",
        16#0ae# => x"ff",
        16#0af# => x"4c",
        16#0b0# => x"98",
        16#0b1# => x"f8",
        16#0b2# => x"a9",
        16#0b3# => x"7e",
        16#0b4# => x"20",
        16#0b5# => x"f4",
        16#0b6# => x"ff",
        16#0b7# => x"00",
        16#0b8# => x"11",
        16#0b9# => x"45",
        16#0ba# => x"73",
        16#0bb# => x"63",
        16#0bc# => x"61",
        16#0bd# => x"70",
        16#0be# => x"65",
        16#0bf# => x"00",
        16#0c0# => x"a5",
        16#0c1# => x"f6",
        16#0c2# => x"85",
        16#0c3# => x"ee",
        16#0c4# => x"85",
        16#0c5# => x"f2",
        16#0c6# => x"a5",
        16#0c7# => x"f7",
        16#0c8# => x"85",
        16#0c9# => x"ef",
        16#0ca# => x"85",
        16#0cb# => x"f3",
        16#0cc# => x"a0",
        16#0cd# => x"07",
        16#0ce# => x"b1",
        16#0cf# => x"ee",
        16#0d0# => x"d8",
        16#0d1# => x"18",
        16#0d2# => x"65",
        16#0d3# => x"ee",
        16#0d4# => x"85",
        16#0d5# => x"fd",
        16#0d6# => x"a9",
        16#0d7# => x"00",
        16#0d8# => x"65",
        16#0d9# => x"ef",
        16#0da# => x"85",
        16#0db# => x"fe",
        16#0dc# => x"a0",
        16#0dd# => x"00",
        16#0de# => x"b1",
        16#0df# => x"fd",
        16#0e0# => x"d0",
        16#0e1# => x"23",
        16#0e2# => x"c8",
        16#0e3# => x"b1",
        16#0e4# => x"fd",
        16#0e5# => x"c9",
        16#0e6# => x"28",
        16#0e7# => x"d0",
        16#0e8# => x"1c",
        16#0e9# => x"c8",
        16#0ea# => x"b1",
        16#0eb# => x"fd",
        16#0ec# => x"c9",
        16#0ed# => x"43",
        16#0ee# => x"d0",
        16#0ef# => x"15",
        16#0f0# => x"c8",
        16#0f1# => x"b1",
        16#0f2# => x"fd",
        16#0f3# => x"c9",
        16#0f4# => x"29",
        16#0f5# => x"d0",
        16#0f6# => x"0e",
        16#0f7# => x"a0",
        16#0f8# => x"06",
        16#0f9# => x"b1",
        16#0fa# => x"ee",
        16#0fb# => x"29",
        16#0fc# => x"4f",
        16#0fd# => x"c9",
        16#0fe# => x"40",
        16#0ff# => x"90",
        16#100# => x"09",
        16#101# => x"29",
        16#102# => x"0d",
        16#103# => x"d0",
        16#104# => x"28",
        16#105# => x"a9",
        16#106# => x"01",
        16#107# => x"6c",
        16#108# => x"f2",
        16#109# => x"00",
        16#10a# => x"a9",
        16#10b# => x"50",
        16#10c# => x"8d",
        16#10d# => x"02",
        16#10e# => x"02",
        16#10f# => x"a9",
        16#110# => x"f9",
        16#111# => x"8d",
        16#112# => x"03",
        16#113# => x"02",
        16#114# => x"00",
        16#115# => x"00",
        16#116# => x"54",
        16#117# => x"68",
        16#118# => x"69",
        16#119# => x"73",
        16#11a# => x"20",
        16#11b# => x"69",
        16#11c# => x"73",
        16#11d# => x"20",
        16#11e# => x"6e",
        16#11f# => x"6f",
        16#120# => x"74",
        16#121# => x"20",
        16#122# => x"61",
        16#123# => x"20",
        16#124# => x"6c",
        16#125# => x"61",
        16#126# => x"6e",
        16#127# => x"67",
        16#128# => x"75",
        16#129# => x"61",
        16#12a# => x"67",
        16#12b# => x"65",
        16#12c# => x"00",
        16#12d# => x"a9",
        16#12e# => x"50",
        16#12f# => x"8d",
        16#130# => x"02",
        16#131# => x"02",
        16#132# => x"a9",
        16#133# => x"f9",
        16#134# => x"8d",
        16#135# => x"03",
        16#136# => x"02",
        16#137# => x"00",
        16#138# => x"00",
        16#139# => x"49",
        16#13a# => x"20",
        16#13b# => x"63",
        16#13c# => x"61",
        16#13d# => x"6e",
        16#13e# => x"6e",
        16#13f# => x"6f",
        16#140# => x"74",
        16#141# => x"20",
        16#142# => x"72",
        16#143# => x"75",
        16#144# => x"6e",
        16#145# => x"20",
        16#146# => x"74",
        16#147# => x"68",
        16#148# => x"69",
        16#149# => x"73",
        16#14a# => x"20",
        16#14b# => x"63",
        16#14c# => x"6f",
        16#14d# => x"64",
        16#14e# => x"65",
        16#14f# => x"00",
        16#150# => x"a2",
        16#151# => x"ff",
        16#152# => x"9a",
        16#153# => x"20",
        16#154# => x"e7",
        16#155# => x"ff",
        16#156# => x"a0",
        16#157# => x"01",
        16#158# => x"b1",
        16#159# => x"fd",
        16#15a# => x"f0",
        16#15b# => x"06",
        16#15c# => x"20",
        16#15d# => x"ee",
        16#15e# => x"ff",
        16#15f# => x"c8",
        16#160# => x"d0",
        16#161# => x"f6",
        16#162# => x"20",
        16#163# => x"e7",
        16#164# => x"ff",
        16#165# => x"4c",
        16#166# => x"98",
        16#167# => x"f8",
        16#168# => x"36",
        16#169# => x"02",
        16#16a# => x"ca",
        16#16b# => x"20",
        16#16c# => x"ff",
        16#16d# => x"2c",
        16#16e# => x"f8",
        16#16f# => x"fe",
        16#170# => x"ea",
        16#171# => x"50",
        16#172# => x"fa",
        16#173# => x"8d",
        16#174# => x"f9",
        16#175# => x"fe",
        16#176# => x"60",
        16#177# => x"a9",
        16#178# => x"00",
        16#179# => x"20",
        16#17a# => x"57",
        16#17b# => x"fc",
        16#17c# => x"20",
        16#17d# => x"80",
        16#17e# => x"f9",
        16#17f# => x"0a",
        16#180# => x"2c",
        16#181# => x"fa",
        16#182# => x"fe",
        16#183# => x"10",
        16#184# => x"fb",
        16#185# => x"ad",
        16#186# => x"fb",
        16#187# => x"fe",
        16#188# => x"60",
        16#189# => x"c8",
        16#18a# => x"b1",
        16#18b# => x"f8",
        16#18c# => x"c9",
        16#18d# => x"20",
        16#18e# => x"f0",
        16#18f# => x"f9",
        16#190# => x"60",
        16#191# => x"a2",
        16#192# => x"00",
        16#193# => x"86",
        16#194# => x"f0",
        16#195# => x"86",
        16#196# => x"f1",
        16#197# => x"b1",
        16#198# => x"f8",
        16#199# => x"c9",
        16#19a# => x"30",
        16#19b# => x"90",
        16#19c# => x"1f",
        16#19d# => x"c9",
        16#19e# => x"3a",
        16#19f# => x"90",
        16#1a0# => x"0a",
        16#1a1# => x"29",
        16#1a2# => x"df",
        16#1a3# => x"e9",
        16#1a4# => x"07",
        16#1a5# => x"90",
        16#1a6# => x"15",
        16#1a7# => x"c9",
        16#1a8# => x"40",
        16#1a9# => x"b0",
        16#1aa# => x"11",
        16#1ab# => x"0a",
        16#1ac# => x"0a",
        16#1ad# => x"0a",
        16#1ae# => x"0a",
        16#1af# => x"a2",
        16#1b0# => x"03",
        16#1b1# => x"0a",
        16#1b2# => x"26",
        16#1b3# => x"f0",
        16#1b4# => x"26",
        16#1b5# => x"f1",
        16#1b6# => x"ca",
        16#1b7# => x"10",
        16#1b8# => x"f8",
        16#1b9# => x"c8",
        16#1ba# => x"d0",
        16#1bb# => x"db",
        16#1bc# => x"60",
        16#1bd# => x"86",
        16#1be# => x"f8",
        16#1bf# => x"84",
        16#1c0# => x"f9",
        16#1c1# => x"a0",
        16#1c2# => x"00",
        16#1c3# => x"2c",
        16#1c4# => x"fa",
        16#1c5# => x"fe",
        16#1c6# => x"50",
        16#1c7# => x"fb",
        16#1c8# => x"b1",
        16#1c9# => x"f8",
        16#1ca# => x"8d",
        16#1cb# => x"fb",
        16#1cc# => x"fe",
        16#1cd# => x"c8",
        16#1ce# => x"c9",
        16#1cf# => x"0d",
        16#1d0# => x"d0",
        16#1d1# => x"f1",
        16#1d2# => x"a4",
        16#1d3# => x"f9",
        16#1d4# => x"60",
        16#1d5# => x"48",
        16#1d6# => x"86",
        16#1d7# => x"f8",
        16#1d8# => x"84",
        16#1d9# => x"f9",
        16#1da# => x"a0",
        16#1db# => x"00",
        16#1dc# => x"20",
        16#1dd# => x"8a",
        16#1de# => x"f9",
        16#1df# => x"c8",
        16#1e0# => x"c9",
        16#1e1# => x"2a",
        16#1e2# => x"f0",
        16#1e3# => x"f8",
        16#1e4# => x"29",
        16#1e5# => x"df",
        16#1e6# => x"aa",
        16#1e7# => x"b1",
        16#1e8# => x"f8",
        16#1e9# => x"e0",
        16#1ea# => x"47",
        16#1eb# => x"f0",
        16#1ec# => x"5e",
        16#1ed# => x"e0",
        16#1ee# => x"48",
        16#1ef# => x"d0",
        16#1f0# => x"49",
        16#1f1# => x"c9",
        16#1f2# => x"2e",
        16#1f3# => x"f0",
        16#1f4# => x"2d",
        16#1f5# => x"29",
        16#1f6# => x"df",
        16#1f7# => x"c9",
        16#1f8# => x"45",
        16#1f9# => x"d0",
        16#1fa# => x"3f",
        16#1fb# => x"c8",
        16#1fc# => x"b1",
        16#1fd# => x"f8",
        16#1fe# => x"c9",
        16#1ff# => x"2e",
        16#200# => x"f0",
        16#201# => x"20",
        16#202# => x"29",
        16#203# => x"df",
        16#204# => x"c9",
        16#205# => x"4c",
        16#206# => x"d0",
        16#207# => x"32",
        16#208# => x"c8",
        16#209# => x"b1",
        16#20a# => x"f8",
        16#20b# => x"c9",
        16#20c# => x"2e",
        16#20d# => x"f0",
        16#20e# => x"13",
        16#20f# => x"29",
        16#210# => x"df",
        16#211# => x"c9",
        16#212# => x"50",
        16#213# => x"d0",
        16#214# => x"25",
        16#215# => x"c8",
        16#216# => x"b1",
        16#217# => x"f8",
        16#218# => x"29",
        16#219# => x"df",
        16#21a# => x"c9",
        16#21b# => x"41",
        16#21c# => x"90",
        16#21d# => x"04",
        16#21e# => x"c9",
        16#21f# => x"5b",
        16#220# => x"90",
        16#221# => x"18",
        16#222# => x"20",
        16#223# => x"a5",
        16#224# => x"fe",
        16#225# => x"0a",
        16#226# => x"0d",
        16#227# => x"36",
        16#228# => x"35",
        16#229# => x"43",
        16#22a# => x"31",
        16#22b# => x"30",
        16#22c# => x"32",
        16#22d# => x"20",
        16#22e# => x"54",
        16#22f# => x"55",
        16#230# => x"42",
        16#231# => x"45",
        16#232# => x"20",
        16#233# => x"31",
        16#234# => x"2e",
        16#235# => x"31",
        16#236# => x"30",
        16#237# => x"0a",
        16#238# => x"0d",
        16#239# => x"ea",
        16#23a# => x"a9",
        16#23b# => x"02",
        16#23c# => x"20",
        16#23d# => x"57",
        16#23e# => x"fc",
        16#23f# => x"20",
        16#240# => x"c1",
        16#241# => x"f9",
        16#242# => x"20",
        16#243# => x"80",
        16#244# => x"f9",
        16#245# => x"c9",
        16#246# => x"80",
        16#247# => x"f0",
        16#248# => x"20",
        16#249# => x"68",
        16#24a# => x"60",
        16#24b# => x"29",
        16#24c# => x"df",
        16#24d# => x"c9",
        16#24e# => x"4f",
        16#24f# => x"d0",
        16#250# => x"e9",
        16#251# => x"20",
        16#252# => x"89",
        16#253# => x"f9",
        16#254# => x"20",
        16#255# => x"91",
        16#256# => x"f9",
        16#257# => x"20",
        16#258# => x"8a",
        16#259# => x"f9",
        16#25a# => x"c9",
        16#25b# => x"0d",
        16#25c# => x"d0",
        16#25d# => x"dc",
        16#25e# => x"8a",
        16#25f# => x"f0",
        16#260# => x"08",
        16#261# => x"a5",
        16#262# => x"f0",
        16#263# => x"85",
        16#264# => x"f6",
        16#265# => x"a5",
        16#266# => x"f1",
        16#267# => x"85",
        16#268# => x"f7",
        16#269# => x"a5",
        16#26a# => x"ef",
        16#26b# => x"48",
        16#26c# => x"a5",
        16#26d# => x"ee",
        16#26e# => x"48",
        16#26f# => x"20",
        16#270# => x"c0",
        16#271# => x"f8",
        16#272# => x"68",
        16#273# => x"85",
        16#274# => x"ee",
        16#275# => x"85",
        16#276# => x"f2",
        16#277# => x"68",
        16#278# => x"85",
        16#279# => x"ef",
        16#27a# => x"85",
        16#27b# => x"f3",
        16#27c# => x"68",
        16#27d# => x"60",
        16#27e# => x"f0",
        16#27f# => x"c2",
        16#280# => x"c9",
        16#281# => x"80",
        16#282# => x"b0",
        16#283# => x"25",
        16#284# => x"48",
        16#285# => x"a9",
        16#286# => x"04",
        16#287# => x"2c",
        16#288# => x"fa",
        16#289# => x"fe",
        16#28a# => x"50",
        16#28b# => x"fb",
        16#28c# => x"8d",
        16#28d# => x"fb",
        16#28e# => x"fe",
        16#28f# => x"2c",
        16#290# => x"fa",
        16#291# => x"fe",
        16#292# => x"50",
        16#293# => x"fb",
        16#294# => x"8e",
        16#295# => x"fb",
        16#296# => x"fe",
        16#297# => x"68",
        16#298# => x"2c",
        16#299# => x"fa",
        16#29a# => x"fe",
        16#29b# => x"50",
        16#29c# => x"fb",
        16#29d# => x"8d",
        16#29e# => x"fb",
        16#29f# => x"fe",
        16#2a0# => x"2c",
        16#2a1# => x"fa",
        16#2a2# => x"fe",
        16#2a3# => x"10",
        16#2a4# => x"fb",
        16#2a5# => x"ae",
        16#2a6# => x"fb",
        16#2a7# => x"fe",
        16#2a8# => x"60",
        16#2a9# => x"c9",
        16#2aa# => x"82",
        16#2ab# => x"f0",
        16#2ac# => x"5a",
        16#2ad# => x"c9",
        16#2ae# => x"83",
        16#2af# => x"f0",
        16#2b0# => x"51",
        16#2b1# => x"c9",
        16#2b2# => x"84",
        16#2b3# => x"f0",
        16#2b4# => x"48",
        16#2b5# => x"48",
        16#2b6# => x"a9",
        16#2b7# => x"06",
        16#2b8# => x"2c",
        16#2b9# => x"fa",
        16#2ba# => x"fe",
        16#2bb# => x"50",
        16#2bc# => x"fb",
        16#2bd# => x"8d",
        16#2be# => x"fb",
        16#2bf# => x"fe",
        16#2c0# => x"2c",
        16#2c1# => x"fa",
        16#2c2# => x"fe",
        16#2c3# => x"50",
        16#2c4# => x"fb",
        16#2c5# => x"8e",
        16#2c6# => x"fb",
        16#2c7# => x"fe",
        16#2c8# => x"2c",
        16#2c9# => x"fa",
        16#2ca# => x"fe",
        16#2cb# => x"50",
        16#2cc# => x"fb",
        16#2cd# => x"8c",
        16#2ce# => x"fb",
        16#2cf# => x"fe",
        16#2d0# => x"68",
        16#2d1# => x"2c",
        16#2d2# => x"fa",
        16#2d3# => x"fe",
        16#2d4# => x"50",
        16#2d5# => x"fb",
        16#2d6# => x"8d",
        16#2d7# => x"fb",
        16#2d8# => x"fe",
        16#2d9# => x"c9",
        16#2da# => x"8e",
        16#2db# => x"f0",
        16#2dc# => x"a1",
        16#2dd# => x"c9",
        16#2de# => x"9d",
        16#2df# => x"f0",
        16#2e0# => x"1b",
        16#2e1# => x"48",
        16#2e2# => x"2c",
        16#2e3# => x"fa",
        16#2e4# => x"fe",
        16#2e5# => x"10",
        16#2e6# => x"fb",
        16#2e7# => x"ad",
        16#2e8# => x"fb",
        16#2e9# => x"fe",
        16#2ea# => x"0a",
        16#2eb# => x"68",
        16#2ec# => x"2c",
        16#2ed# => x"fa",
        16#2ee# => x"fe",
        16#2ef# => x"10",
        16#2f0# => x"fb",
        16#2f1# => x"ac",
        16#2f2# => x"fb",
        16#2f3# => x"fe",
        16#2f4# => x"2c",
        16#2f5# => x"fa",
        16#2f6# => x"fe",
        16#2f7# => x"10",
        16#2f8# => x"fb",
        16#2f9# => x"ae",
        16#2fa# => x"fb",
        16#2fb# => x"fe",
        16#2fc# => x"60",
        16#2fd# => x"a6",
        16#2fe# => x"f2",
        16#2ff# => x"a4",
        16#300# => x"f3",
        16#301# => x"60",
        16#302# => x"a2",
        16#303# => x"00",
        16#304# => x"a0",
        16#305# => x"08",
        16#306# => x"60",
        16#307# => x"a2",
        16#308# => x"00",
        16#309# => x"a0",
        16#30a# => x"00",
        16#30b# => x"60",
        16#30c# => x"86",
        16#30d# => x"f8",
        16#30e# => x"84",
        16#30f# => x"f9",
        16#310# => x"a8",
        16#311# => x"f0",
        16#312# => x"71",
        16#313# => x"48",
        16#314# => x"a0",
        16#315# => x"08",
        16#316# => x"2c",
        16#317# => x"fa",
        16#318# => x"fe",
        16#319# => x"50",
        16#31a# => x"fb",
        16#31b# => x"8c",
        16#31c# => x"fb",
        16#31d# => x"fe",
        16#31e# => x"2c",
        16#31f# => x"fa",
        16#320# => x"fe",
        16#321# => x"50",
        16#322# => x"fb",
        16#323# => x"8d",
        16#324# => x"fb",
        16#325# => x"fe",
        16#326# => x"aa",
        16#327# => x"10",
        16#328# => x"08",
        16#329# => x"a0",
        16#32a# => x"00",
        16#32b# => x"b1",
        16#32c# => x"f8",
        16#32d# => x"a8",
        16#32e# => x"4c",
        16#32f# => x"3a",
        16#330# => x"fb",
        16#331# => x"bc",
        16#332# => x"c9",
        16#333# => x"fc",
        16#334# => x"e0",
        16#335# => x"15",
        16#336# => x"90",
        16#337# => x"02",
        16#338# => x"a0",
        16#339# => x"10",
        16#33a# => x"2c",
        16#33b# => x"fa",
        16#33c# => x"fe",
        16#33d# => x"50",
        16#33e# => x"fb",
        16#33f# => x"8c",
        16#340# => x"fb",
        16#341# => x"fe",
        16#342# => x"88",
        16#343# => x"30",
        16#344# => x"0d",
        16#345# => x"2c",
        16#346# => x"fa",
        16#347# => x"fe",
        16#348# => x"50",
        16#349# => x"fb",
        16#34a# => x"b1",
        16#34b# => x"f8",
        16#34c# => x"8d",
        16#34d# => x"fb",
        16#34e# => x"fe",
        16#34f# => x"88",
        16#350# => x"10",
        16#351# => x"f3",
        16#352# => x"8a",
        16#353# => x"10",
        16#354# => x"08",
        16#355# => x"a0",
        16#356# => x"01",
        16#357# => x"b1",
        16#358# => x"f8",
        16#359# => x"a8",
        16#35a# => x"4c",
        16#35b# => x"66",
        16#35c# => x"fb",
        16#35d# => x"bc",
        16#35e# => x"dd",
        16#35f# => x"fc",
        16#360# => x"e0",
        16#361# => x"15",
        16#362# => x"90",
        16#363# => x"02",
        16#364# => x"a0",
        16#365# => x"10",
        16#366# => x"2c",
        16#367# => x"fa",
        16#368# => x"fe",
        16#369# => x"50",
        16#36a# => x"fb",
        16#36b# => x"8c",
        16#36c# => x"fb",
        16#36d# => x"fe",
        16#36e# => x"88",
        16#36f# => x"30",
        16#370# => x"0d",
        16#371# => x"2c",
        16#372# => x"fa",
        16#373# => x"fe",
        16#374# => x"10",
        16#375# => x"fb",
        16#376# => x"ad",
        16#377# => x"fb",
        16#378# => x"fe",
        16#379# => x"91",
        16#37a# => x"f8",
        16#37b# => x"88",
        16#37c# => x"10",
        16#37d# => x"f3",
        16#37e# => x"a4",
        16#37f# => x"f9",
        16#380# => x"a6",
        16#381# => x"f8",
        16#382# => x"68",
        16#383# => x"60",
        16#384# => x"a9",
        16#385# => x"0a",
        16#386# => x"20",
        16#387# => x"57",
        16#388# => x"fc",
        16#389# => x"a0",
        16#38a# => x"04",
        16#38b# => x"2c",
        16#38c# => x"fa",
        16#38d# => x"fe",
        16#38e# => x"50",
        16#38f# => x"fb",
        16#390# => x"b1",
        16#391# => x"f8",
        16#392# => x"8d",
        16#393# => x"fb",
        16#394# => x"fe",
        16#395# => x"88",
        16#396# => x"c0",
        16#397# => x"01",
        16#398# => x"d0",
        16#399# => x"f1",
        16#39a# => x"a9",
        16#39b# => x"07",
        16#39c# => x"20",
        16#39d# => x"57",
        16#39e# => x"fc",
        16#39f# => x"b1",
        16#3a0# => x"f8",
        16#3a1# => x"48",
        16#3a2# => x"88",
        16#3a3# => x"2c",
        16#3a4# => x"fa",
        16#3a5# => x"fe",
        16#3a6# => x"50",
        16#3a7# => x"fb",
        16#3a8# => x"8c",
        16#3a9# => x"fb",
        16#3aa# => x"fe",
        16#3ab# => x"b1",
        16#3ac# => x"f8",
        16#3ad# => x"48",
        16#3ae# => x"a2",
        16#3af# => x"ff",
        16#3b0# => x"20",
        16#3b1# => x"80",
        16#3b2# => x"f9",
        16#3b3# => x"c9",
        16#3b4# => x"80",
        16#3b5# => x"b0",
        16#3b6# => x"1d",
        16#3b7# => x"68",
        16#3b8# => x"85",
        16#3b9# => x"f8",
        16#3ba# => x"68",
        16#3bb# => x"85",
        16#3bc# => x"f9",
        16#3bd# => x"a0",
        16#3be# => x"00",
        16#3bf# => x"2c",
        16#3c0# => x"fa",
        16#3c1# => x"fe",
        16#3c2# => x"10",
        16#3c3# => x"fb",
        16#3c4# => x"ad",
        16#3c5# => x"fb",
        16#3c6# => x"fe",
        16#3c7# => x"91",
        16#3c8# => x"f8",
        16#3c9# => x"c8",
        16#3ca# => x"c9",
        16#3cb# => x"0d",
        16#3cc# => x"d0",
        16#3cd# => x"f1",
        16#3ce# => x"a9",
        16#3cf# => x"00",
        16#3d0# => x"88",
        16#3d1# => x"18",
        16#3d2# => x"e8",
        16#3d3# => x"60",
        16#3d4# => x"68",
        16#3d5# => x"68",
        16#3d6# => x"a9",
        16#3d7# => x"00",
        16#3d8# => x"60",
        16#3d9# => x"48",
        16#3da# => x"a9",
        16#3db# => x"0c",
        16#3dc# => x"20",
        16#3dd# => x"57",
        16#3de# => x"fc",
        16#3df# => x"2c",
        16#3e0# => x"fa",
        16#3e1# => x"fe",
        16#3e2# => x"50",
        16#3e3# => x"fb",
        16#3e4# => x"8c",
        16#3e5# => x"fb",
        16#3e6# => x"fe",
        16#3e7# => x"b5",
        16#3e8# => x"03",
        16#3e9# => x"20",
        16#3ea# => x"57",
        16#3eb# => x"fc",
        16#3ec# => x"b5",
        16#3ed# => x"02",
        16#3ee# => x"20",
        16#3ef# => x"57",
        16#3f0# => x"fc",
        16#3f1# => x"b5",
        16#3f2# => x"01",
        16#3f3# => x"20",
        16#3f4# => x"57",
        16#3f5# => x"fc",
        16#3f6# => x"b5",
        16#3f7# => x"00",
        16#3f8# => x"20",
        16#3f9# => x"57",
        16#3fa# => x"fc",
        16#3fb# => x"68",
        16#3fc# => x"20",
        16#3fd# => x"57",
        16#3fe# => x"fc",
        16#3ff# => x"20",
        16#400# => x"80",
        16#401# => x"f9",
        16#402# => x"48",
        16#403# => x"20",
        16#404# => x"80",
        16#405# => x"f9",
        16#406# => x"95",
        16#407# => x"03",
        16#408# => x"20",
        16#409# => x"80",
        16#40a# => x"f9",
        16#40b# => x"95",
        16#40c# => x"02",
        16#40d# => x"20",
        16#40e# => x"80",
        16#40f# => x"f9",
        16#410# => x"95",
        16#411# => x"01",
        16#412# => x"20",
        16#413# => x"80",
        16#414# => x"f9",
        16#415# => x"95",
        16#416# => x"00",
        16#417# => x"68",
        16#418# => x"60",
        16#419# => x"48",
        16#41a# => x"a9",
        16#41b# => x"12",
        16#41c# => x"20",
        16#41d# => x"57",
        16#41e# => x"fc",
        16#41f# => x"68",
        16#420# => x"20",
        16#421# => x"57",
        16#422# => x"fc",
        16#423# => x"c9",
        16#424# => x"00",
        16#425# => x"d0",
        16#426# => x"0a",
        16#427# => x"48",
        16#428# => x"98",
        16#429# => x"20",
        16#42a# => x"57",
        16#42b# => x"fc",
        16#42c# => x"20",
        16#42d# => x"80",
        16#42e# => x"f9",
        16#42f# => x"68",
        16#430# => x"60",
        16#431# => x"20",
        16#432# => x"bd",
        16#433# => x"f9",
        16#434# => x"4c",
        16#435# => x"80",
        16#436# => x"f9",
        16#437# => x"a9",
        16#438# => x"0e",
        16#439# => x"20",
        16#43a# => x"57",
        16#43b# => x"fc",
        16#43c# => x"98",
        16#43d# => x"20",
        16#43e# => x"57",
        16#43f# => x"fc",
        16#440# => x"4c",
        16#441# => x"7c",
        16#442# => x"f9",
        16#443# => x"48",
        16#444# => x"a9",
        16#445# => x"10",
        16#446# => x"20",
        16#447# => x"57",
        16#448# => x"fc",
        16#449# => x"98",
        16#44a# => x"20",
        16#44b# => x"57",
        16#44c# => x"fc",
        16#44d# => x"68",
        16#44e# => x"20",
        16#44f# => x"57",
        16#450# => x"fc",
        16#451# => x"48",
        16#452# => x"20",
        16#453# => x"80",
        16#454# => x"f9",
        16#455# => x"68",
        16#456# => x"60",
        16#457# => x"2c",
        16#458# => x"fa",
        16#459# => x"fe",
        16#45a# => x"50",
        16#45b# => x"fb",
        16#45c# => x"8d",
        16#45d# => x"fb",
        16#45e# => x"fe",
        16#45f# => x"60",
        16#460# => x"84",
        16#461# => x"fb",
        16#462# => x"86",
        16#463# => x"fa",
        16#464# => x"48",
        16#465# => x"a9",
        16#466# => x"14",
        16#467# => x"20",
        16#468# => x"57",
        16#469# => x"fc",
        16#46a# => x"a0",
        16#46b# => x"11",
        16#46c# => x"b1",
        16#46d# => x"fa",
        16#46e# => x"20",
        16#46f# => x"57",
        16#470# => x"fc",
        16#471# => x"88",
        16#472# => x"c0",
        16#473# => x"01",
        16#474# => x"d0",
        16#475# => x"f6",
        16#476# => x"88",
        16#477# => x"b1",
        16#478# => x"fa",
        16#479# => x"aa",
        16#47a# => x"c8",
        16#47b# => x"b1",
        16#47c# => x"fa",
        16#47d# => x"a8",
        16#47e# => x"20",
        16#47f# => x"bd",
        16#480# => x"f9",
        16#481# => x"68",
        16#482# => x"20",
        16#483# => x"57",
        16#484# => x"fc",
        16#485# => x"20",
        16#486# => x"80",
        16#487# => x"f9",
        16#488# => x"48",
        16#489# => x"a0",
        16#48a# => x"11",
        16#48b# => x"20",
        16#48c# => x"80",
        16#48d# => x"f9",
        16#48e# => x"91",
        16#48f# => x"fa",
        16#490# => x"88",
        16#491# => x"c0",
        16#492# => x"01",
        16#493# => x"d0",
        16#494# => x"f6",
        16#495# => x"a4",
        16#496# => x"fb",
        16#497# => x"a6",
        16#498# => x"fa",
        16#499# => x"68",
        16#49a# => x"60",
        16#49b# => x"84",
        16#49c# => x"fb",
        16#49d# => x"86",
        16#49e# => x"fa",
        16#49f# => x"48",
        16#4a0# => x"a9",
        16#4a1# => x"16",
        16#4a2# => x"20",
        16#4a3# => x"57",
        16#4a4# => x"fc",
        16#4a5# => x"a0",
        16#4a6# => x"0c",
        16#4a7# => x"b1",
        16#4a8# => x"fa",
        16#4a9# => x"20",
        16#4aa# => x"57",
        16#4ab# => x"fc",
        16#4ac# => x"88",
        16#4ad# => x"10",
        16#4ae# => x"f8",
        16#4af# => x"68",
        16#4b0# => x"20",
        16#4b1# => x"57",
        16#4b2# => x"fc",
        16#4b3# => x"a0",
        16#4b4# => x"0c",
        16#4b5# => x"20",
        16#4b6# => x"80",
        16#4b7# => x"f9",
        16#4b8# => x"91",
        16#4b9# => x"fa",
        16#4ba# => x"88",
        16#4bb# => x"10",
        16#4bc# => x"f8",
        16#4bd# => x"a4",
        16#4be# => x"fb",
        16#4bf# => x"a6",
        16#4c0# => x"fa",
        16#4c1# => x"4c",
        16#4c2# => x"7c",
        16#4c3# => x"f9",
        16#4c4# => x"00",
        16#4c5# => x"ff",
        16#4c6# => x"42",
        16#4c7# => x"61",
        16#4c8# => x"64",
        16#4c9# => x"00",
        16#4ca# => x"00",
        16#4cb# => x"05",
        16#4cc# => x"00",
        16#4cd# => x"05",
        16#4ce# => x"04",
        16#4cf# => x"05",
        16#4d0# => x"08",
        16#4d1# => x"0e",
        16#4d2# => x"04",
        16#4d3# => x"01",
        16#4d4# => x"01",
        16#4d5# => x"05",
        16#4d6# => x"00",
        16#4d7# => x"01",
        16#4d8# => x"20",
        16#4d9# => x"10",
        16#4da# => x"0d",
        16#4db# => x"00",
        16#4dc# => x"04",
        16#4dd# => x"80",
        16#4de# => x"05",
        16#4df# => x"00",
        16#4e0# => x"05",
        16#4e1# => x"00",
        16#4e2# => x"05",
        16#4e3# => x"00",
        16#4e4# => x"00",
        16#4e5# => x"00",
        16#4e6# => x"05",
        16#4e7# => x"09",
        16#4e8# => x"05",
        16#4e9# => x"00",
        16#4ea# => x"08",
        16#4eb# => x"18",
        16#4ec# => x"00",
        16#4ed# => x"01",
        16#4ee# => x"0d",
        16#4ef# => x"80",
        16#4f0# => x"04",
        16#4f1# => x"80",
        16#4f2# => x"85",
        16#4f3# => x"fc",
        16#4f4# => x"68",
        16#4f5# => x"48",
        16#4f6# => x"29",
        16#4f7# => x"10",
        16#4f8# => x"d0",
        16#4f9# => x"10",
        16#4fa# => x"6c",
        16#4fb# => x"04",
        16#4fc# => x"02",
        16#4fd# => x"2c",
        16#4fe# => x"fe",
        16#4ff# => x"fe",
        16#500# => x"30",
        16#501# => x"4a",
        16#502# => x"2c",
        16#503# => x"f8",
        16#504# => x"fe",
        16#505# => x"30",
        16#506# => x"1e",
        16#507# => x"6c",
        16#508# => x"06",
        16#509# => x"02",
        16#50a# => x"8a",
        16#50b# => x"48",
        16#50c# => x"ba",
        16#50d# => x"bd",
        16#50e# => x"03",
        16#50f# => x"01",
        16#510# => x"d8",
        16#511# => x"38",
        16#512# => x"e9",
        16#513# => x"01",
        16#514# => x"85",
        16#515# => x"fd",
        16#516# => x"bd",
        16#517# => x"04",
        16#518# => x"01",
        16#519# => x"e9",
        16#51a# => x"00",
        16#51b# => x"85",
        16#51c# => x"fe",
        16#51d# => x"68",
        16#51e# => x"aa",
        16#51f# => x"a5",
        16#520# => x"fc",
        16#521# => x"58",
        16#522# => x"6c",
        16#523# => x"02",
        16#524# => x"02",
        16#525# => x"ad",
        16#526# => x"f9",
        16#527# => x"fe",
        16#528# => x"30",
        16#529# => x"1c",
        16#52a# => x"98",
        16#52b# => x"48",
        16#52c# => x"8a",
        16#52d# => x"48",
        16#52e# => x"20",
        16#52f# => x"8d",
        16#530# => x"fe",
        16#531# => x"a8",
        16#532# => x"20",
        16#533# => x"8d",
        16#534# => x"fe",
        16#535# => x"aa",
        16#536# => x"20",
        16#537# => x"8d",
        16#538# => x"fe",
        16#539# => x"20",
        16#53a# => x"43",
        16#53b# => x"fd",
        16#53c# => x"68",
        16#53d# => x"aa",
        16#53e# => x"68",
        16#53f# => x"a8",
        16#540# => x"a5",
        16#541# => x"fc",
        16#542# => x"40",
        16#543# => x"6c",
        16#544# => x"20",
        16#545# => x"02",
        16#546# => x"0a",
        16#547# => x"85",
        16#548# => x"ff",
        16#549# => x"a5",
        16#54a# => x"fc",
        16#54b# => x"40",
        16#54c# => x"ad",
        16#54d# => x"ff",
        16#54e# => x"fe",
        16#54f# => x"10",
        16#550# => x"21",
        16#551# => x"58",
        16#552# => x"2c",
        16#553# => x"fa",
        16#554# => x"fe",
        16#555# => x"10",
        16#556# => x"fb",
        16#557# => x"ad",
        16#558# => x"fb",
        16#559# => x"fe",
        16#55a# => x"a9",
        16#55b# => x"00",
        16#55c# => x"8d",
        16#55d# => x"36",
        16#55e# => x"02",
        16#55f# => x"a8",
        16#560# => x"20",
        16#561# => x"80",
        16#562# => x"f9",
        16#563# => x"8d",
        16#564# => x"37",
        16#565# => x"02",
        16#566# => x"c8",
        16#567# => x"20",
        16#568# => x"80",
        16#569# => x"f9",
        16#56a# => x"99",
        16#56b# => x"37",
        16#56c# => x"02",
        16#56d# => x"d0",
        16#56e# => x"f7",
        16#56f# => x"4c",
        16#570# => x"36",
        16#571# => x"02",
        16#572# => x"8d",
        16#573# => x"fa",
        16#574# => x"ff",
        16#575# => x"98",
        16#576# => x"48",
        16#577# => x"ac",
        16#578# => x"fa",
        16#579# => x"ff",
        16#57a# => x"b9",
        16#57b# => x"7d",
        16#57c# => x"fe",
        16#57d# => x"8d",
        16#57e# => x"fa",
        16#57f# => x"ff",
        16#580# => x"b9",
        16#581# => x"85",
        16#582# => x"fe",
        16#583# => x"8d",
        16#584# => x"fb",
        16#585# => x"ff",
        16#586# => x"b9",
        16#587# => x"6d",
        16#588# => x"fe",
        16#589# => x"85",
        16#58a# => x"f4",
        16#58b# => x"b9",
        16#58c# => x"75",
        16#58d# => x"fe",
        16#58e# => x"85",
        16#58f# => x"f5",
        16#590# => x"2c",
        16#591# => x"fe",
        16#592# => x"fe",
        16#593# => x"10",
        16#594# => x"fb",
        16#595# => x"ad",
        16#596# => x"ff",
        16#597# => x"fe",
        16#598# => x"c0",
        16#599# => x"05",
        16#59a# => x"f0",
        16#59b# => x"58",
        16#59c# => x"98",
        16#59d# => x"48",
        16#59e# => x"a0",
        16#59f# => x"01",
        16#5a0# => x"2c",
        16#5a1# => x"fe",
        16#5a2# => x"fe",
        16#5a3# => x"10",
        16#5a4# => x"fb",
        16#5a5# => x"ad",
        16#5a6# => x"ff",
        16#5a7# => x"fe",
        16#5a8# => x"2c",
        16#5a9# => x"fe",
        16#5aa# => x"fe",
        16#5ab# => x"10",
        16#5ac# => x"fb",
        16#5ad# => x"ad",
        16#5ae# => x"ff",
        16#5af# => x"fe",
        16#5b0# => x"2c",
        16#5b1# => x"fe",
        16#5b2# => x"fe",
        16#5b3# => x"10",
        16#5b4# => x"fb",
        16#5b5# => x"ad",
        16#5b6# => x"ff",
        16#5b7# => x"fe",
        16#5b8# => x"91",
        16#5b9# => x"f4",
        16#5ba# => x"88",
        16#5bb# => x"2c",
        16#5bc# => x"fe",
        16#5bd# => x"fe",
        16#5be# => x"10",
        16#5bf# => x"fb",
        16#5c0# => x"ad",
        16#5c1# => x"ff",
        16#5c2# => x"fe",
        16#5c3# => x"91",
        16#5c4# => x"f4",
        16#5c5# => x"2c",
        16#5c6# => x"fd",
        16#5c7# => x"fe",
        16#5c8# => x"2c",
        16#5c9# => x"fd",
        16#5ca# => x"fe",
        16#5cb# => x"2c",
        16#5cc# => x"fe",
        16#5cd# => x"fe",
        16#5ce# => x"10",
        16#5cf# => x"fb",
        16#5d0# => x"ad",
        16#5d1# => x"ff",
        16#5d2# => x"fe",
        16#5d3# => x"68",
        16#5d4# => x"c9",
        16#5d5# => x"06",
        16#5d6# => x"90",
        16#5d7# => x"1c",
        16#5d8# => x"d0",
        16#5d9# => x"1f",
        16#5da# => x"a0",
        16#5db# => x"00",
        16#5dc# => x"ad",
        16#5dd# => x"fc",
        16#5de# => x"fe",
        16#5df# => x"29",
        16#5e0# => x"80",
        16#5e1# => x"10",
        16#5e2# => x"f9",
        16#5e3# => x"b9",
        16#5e4# => x"ff",
        16#5e5# => x"ff",
        16#5e6# => x"8d",
        16#5e7# => x"fd",
        16#5e8# => x"fe",
        16#5e9# => x"c8",
        16#5ea# => x"d0",
        16#5eb# => x"f0",
        16#5ec# => x"2c",
        16#5ed# => x"fc",
        16#5ee# => x"fe",
        16#5ef# => x"10",
        16#5f0# => x"fb",
        16#5f1# => x"8d",
        16#5f2# => x"fd",
        16#5f3# => x"fe",
        16#5f4# => x"68",
        16#5f5# => x"a8",
        16#5f6# => x"a5",
        16#5f7# => x"fc",
        16#5f8# => x"40",
        16#5f9# => x"a0",
        16#5fa# => x"00",
        16#5fb# => x"ad",
        16#5fc# => x"fc",
        16#5fd# => x"fe",
        16#5fe# => x"29",
        16#5ff# => x"80",
        16#600# => x"10",
        16#601# => x"f9",
        16#602# => x"ad",
        16#603# => x"fd",
        16#604# => x"fe",
        16#605# => x"99",
        16#606# => x"ff",
        16#607# => x"ff",
        16#608# => x"c8",
        16#609# => x"d0",
        16#60a# => x"f0",
        16#60b# => x"f0",
        16#60c# => x"e7",
        16#60d# => x"48",
        16#60e# => x"ad",
        16#60f# => x"ff",
        16#610# => x"ff",
        16#611# => x"8d",
        16#612# => x"fd",
        16#613# => x"fe",
        16#614# => x"ee",
        16#615# => x"0f",
        16#616# => x"fe",
        16#617# => x"d0",
        16#618# => x"03",
        16#619# => x"ee",
        16#61a# => x"10",
        16#61b# => x"fe",
        16#61c# => x"68",
        16#61d# => x"40",
        16#61e# => x"48",
        16#61f# => x"ad",
        16#620# => x"fd",
        16#621# => x"fe",
        16#622# => x"8d",
        16#623# => x"ff",
        16#624# => x"ff",
        16#625# => x"ee",
        16#626# => x"23",
        16#627# => x"fe",
        16#628# => x"d0",
        16#629# => x"03",
        16#62a# => x"ee",
        16#62b# => x"24",
        16#62c# => x"fe",
        16#62d# => x"68",
        16#62e# => x"40",
        16#62f# => x"48",
        16#630# => x"98",
        16#631# => x"48",
        16#632# => x"a0",
        16#633# => x"00",
        16#634# => x"b1",
        16#635# => x"f6",
        16#636# => x"8d",
        16#637# => x"fd",
        16#638# => x"fe",
        16#639# => x"e6",
        16#63a# => x"f6",
        16#63b# => x"d0",
        16#63c# => x"02",
        16#63d# => x"e6",
        16#63e# => x"f7",
        16#63f# => x"b1",
        16#640# => x"f6",
        16#641# => x"8d",
        16#642# => x"fd",
        16#643# => x"fe",
        16#644# => x"e6",
        16#645# => x"f6",
        16#646# => x"d0",
        16#647# => x"02",
        16#648# => x"e6",
        16#649# => x"f7",
        16#64a# => x"68",
        16#64b# => x"a8",
        16#64c# => x"68",
        16#64d# => x"40",
        16#64e# => x"48",
        16#64f# => x"98",
        16#650# => x"48",
        16#651# => x"a0",
        16#652# => x"00",
        16#653# => x"ad",
        16#654# => x"fd",
        16#655# => x"fe",
        16#656# => x"91",
        16#657# => x"f6",
        16#658# => x"e6",
        16#659# => x"f6",
        16#65a# => x"d0",
        16#65b# => x"02",
        16#65c# => x"e6",
        16#65d# => x"f7",
        16#65e# => x"ad",
        16#65f# => x"fd",
        16#660# => x"fe",
        16#661# => x"91",
        16#662# => x"f6",
        16#663# => x"e6",
        16#664# => x"f6",
        16#665# => x"d0",
        16#666# => x"02",
        16#667# => x"e6",
        16#668# => x"f7",
        16#669# => x"68",
        16#66a# => x"a8",
        16#66b# => x"68",
        16#66c# => x"40",
        16#66d# => x"0f",
        16#66e# => x"23",
        16#66f# => x"f6",
        16#670# => x"f6",
        16#671# => x"f6",
        16#672# => x"f6",
        16#673# => x"e4",
        16#674# => x"06",
        16#675# => x"fe",
        16#676# => x"fe",
        16#677# => x"00",
        16#678# => x"00",
        16#679# => x"00",
        16#67a# => x"00",
        16#67b# => x"fd",
        16#67c# => x"fe",
        16#67d# => x"0d",
        16#67e# => x"1e",
        16#67f# => x"2f",
        16#680# => x"4e",
        16#681# => x"c0",
        16#682# => x"c0",
        16#683# => x"c0",
        16#684# => x"c0",
        16#685# => x"fe",
        16#686# => x"fe",
        16#687# => x"fe",
        16#688# => x"fe",
        16#689# => x"fe",
        16#68a# => x"fe",
        16#68b# => x"fe",
        16#68c# => x"fe",
        16#68d# => x"2c",
        16#68e# => x"f8",
        16#68f# => x"fe",
        16#690# => x"30",
        16#691# => x"0f",
        16#692# => x"2c",
        16#693# => x"fe",
        16#694# => x"fe",
        16#695# => x"10",
        16#696# => x"f6",
        16#697# => x"a5",
        16#698# => x"fc",
        16#699# => x"08",
        16#69a# => x"58",
        16#69b# => x"28",
        16#69c# => x"85",
        16#69d# => x"fc",
        16#69e# => x"4c",
        16#69f# => x"8d",
        16#6a0# => x"fe",
        16#6a1# => x"ad",
        16#6a2# => x"f9",
        16#6a3# => x"fe",
        16#6a4# => x"60",
        16#6a5# => x"68",
        16#6a6# => x"85",
        16#6a7# => x"fa",
        16#6a8# => x"68",
        16#6a9# => x"85",
        16#6aa# => x"fb",
        16#6ab# => x"a0",
        16#6ac# => x"00",
        16#6ad# => x"e6",
        16#6ae# => x"fa",
        16#6af# => x"d0",
        16#6b0# => x"02",
        16#6b1# => x"e6",
        16#6b2# => x"fb",
        16#6b3# => x"b1",
        16#6b4# => x"fa",
        16#6b5# => x"30",
        16#6b6# => x"06",
        16#6b7# => x"20",
        16#6b8# => x"ee",
        16#6b9# => x"ff",
        16#6ba# => x"4c",
        16#6bb# => x"ad",
        16#6bc# => x"fe",
        16#6bd# => x"6c",
        16#6be# => x"fa",
        16#6bf# => x"00",
        16#6c0# => x"8d",
        16#6c1# => x"fd",
        16#6c2# => x"fe",
        16#6c3# => x"40",
        16#6c4# => x"ff",
        16#6c5# => x"ff",
        16#6c6# => x"ff",
        16#6c7# => x"ff",
        16#6c8# => x"ff",
        16#6c9# => x"ff",
        16#6ca# => x"ff",
        16#6cb# => x"ff",
        16#6cc# => x"ff",
        16#6cd# => x"ff",
        16#6ce# => x"ff",
        16#6cf# => x"ff",
        16#6d0# => x"ff",
        16#6d1# => x"ff",
        16#6d2# => x"ff",
        16#6d3# => x"ff",
        16#6d4# => x"ff",
        16#6d5# => x"ff",
        16#6d6# => x"ff",
        16#6d7# => x"ff",
        16#6d8# => x"ff",
        16#6d9# => x"ff",
        16#6da# => x"ff",
        16#6db# => x"ff",
        16#6dc# => x"ff",
        16#6dd# => x"ff",
        16#6de# => x"ff",
        16#6df# => x"ff",
        16#6e0# => x"ff",
        16#6e1# => x"ff",
        16#6e2# => x"ff",
        16#6e3# => x"ff",
        16#6e4# => x"ff",
        16#6e5# => x"ff",
        16#6e6# => x"ff",
        16#6e7# => x"ff",
        16#6e8# => x"ff",
        16#6e9# => x"ff",
        16#6ea# => x"ff",
        16#6eb# => x"ff",
        16#6ec# => x"ff",
        16#6ed# => x"ff",
        16#6ee# => x"ff",
        16#6ef# => x"ff",
        16#6f0# => x"00",
        16#6f1# => x"00",
        16#6f2# => x"00",
        16#6f3# => x"00",
        16#6f4# => x"00",
        16#6f5# => x"00",
        16#6f6# => x"00",
        16#6f7# => x"00",
        16#6f8# => x"00",
        16#6f9# => x"00",
        16#6fa# => x"00",
        16#6fb# => x"00",
        16#6fc# => x"00",
        16#6fd# => x"00",
        16#6fe# => x"00",
        16#6ff# => x"00",
        16#700# => x"ff",
        16#701# => x"ff",
        16#702# => x"ff",
        16#703# => x"ff",
        16#704# => x"ff",
        16#705# => x"ff",
        16#706# => x"ff",
        16#707# => x"ff",
        16#708# => x"ff",
        16#709# => x"ff",
        16#70a# => x"ff",
        16#70b# => x"ff",
        16#70c# => x"ff",
        16#70d# => x"ff",
        16#70e# => x"ff",
        16#70f# => x"ff",
        16#710# => x"ff",
        16#711# => x"ff",
        16#712# => x"ff",
        16#713# => x"ff",
        16#714# => x"ff",
        16#715# => x"ff",
        16#716# => x"ff",
        16#717# => x"ff",
        16#718# => x"ff",
        16#719# => x"ff",
        16#71a# => x"ff",
        16#71b# => x"ff",
        16#71c# => x"ff",
        16#71d# => x"ff",
        16#71e# => x"ff",
        16#71f# => x"ff",
        16#720# => x"ff",
        16#721# => x"ff",
        16#722# => x"ff",
        16#723# => x"ff",
        16#724# => x"ff",
        16#725# => x"ff",
        16#726# => x"ff",
        16#727# => x"ff",
        16#728# => x"ff",
        16#729# => x"ff",
        16#72a# => x"ff",
        16#72b# => x"ff",
        16#72c# => x"ff",
        16#72d# => x"ff",
        16#72e# => x"ff",
        16#72f# => x"ff",
        16#730# => x"ff",
        16#731# => x"ff",
        16#732# => x"ff",
        16#733# => x"ff",
        16#734# => x"ff",
        16#735# => x"ff",
        16#736# => x"ff",
        16#737# => x"ff",
        16#738# => x"ff",
        16#739# => x"ff",
        16#73a# => x"ff",
        16#73b# => x"ff",
        16#73c# => x"ff",
        16#73d# => x"ff",
        16#73e# => x"ff",
        16#73f# => x"ff",
        16#740# => x"ff",
        16#741# => x"ff",
        16#742# => x"ff",
        16#743# => x"ff",
        16#744# => x"ff",
        16#745# => x"ff",
        16#746# => x"ff",
        16#747# => x"ff",
        16#748# => x"ff",
        16#749# => x"ff",
        16#74a# => x"ff",
        16#74b# => x"ff",
        16#74c# => x"ff",
        16#74d# => x"ff",
        16#74e# => x"ff",
        16#74f# => x"ff",
        16#750# => x"ff",
        16#751# => x"ff",
        16#752# => x"ff",
        16#753# => x"ff",
        16#754# => x"ff",
        16#755# => x"ff",
        16#756# => x"ff",
        16#757# => x"ff",
        16#758# => x"ff",
        16#759# => x"ff",
        16#75a# => x"ff",
        16#75b# => x"ff",
        16#75c# => x"ff",
        16#75d# => x"ff",
        16#75e# => x"ff",
        16#75f# => x"ff",
        16#760# => x"ff",
        16#761# => x"ff",
        16#762# => x"ff",
        16#763# => x"ff",
        16#764# => x"ff",
        16#765# => x"ff",
        16#766# => x"ff",
        16#767# => x"ff",
        16#768# => x"ff",
        16#769# => x"ff",
        16#76a# => x"ff",
        16#76b# => x"ff",
        16#76c# => x"ff",
        16#76d# => x"ff",
        16#76e# => x"ff",
        16#76f# => x"ff",
        16#770# => x"ff",
        16#771# => x"ff",
        16#772# => x"ff",
        16#773# => x"ff",
        16#774# => x"ff",
        16#775# => x"ff",
        16#776# => x"ff",
        16#777# => x"ff",
        16#778# => x"ff",
        16#779# => x"ff",
        16#77a# => x"ff",
        16#77b# => x"ff",
        16#77c# => x"ff",
        16#77d# => x"ff",
        16#77e# => x"ff",
        16#77f# => x"ff",
        16#780# => x"c4",
        16#781# => x"fc",
        16#782# => x"50",
        16#783# => x"f9",
        16#784# => x"fd",
        16#785# => x"fc",
        16#786# => x"c4",
        16#787# => x"fc",
        16#788# => x"d5",
        16#789# => x"f9",
        16#78a# => x"80",
        16#78b# => x"fa",
        16#78c# => x"0c",
        16#78d# => x"fb",
        16#78e# => x"6d",
        16#78f# => x"f9",
        16#790# => x"77",
        16#791# => x"f9",
        16#792# => x"60",
        16#793# => x"fc",
        16#794# => x"d9",
        16#795# => x"fb",
        16#796# => x"37",
        16#797# => x"fc",
        16#798# => x"43",
        16#799# => x"fc",
        16#79a# => x"9b",
        16#79b# => x"fc",
        16#79c# => x"19",
        16#79d# => x"fc",
        16#79e# => x"c4",
        16#79f# => x"fc",
        16#7a0# => x"88",
        16#7a1# => x"f9",
        16#7a2# => x"c4",
        16#7a3# => x"fc",
        16#7a4# => x"c4",
        16#7a5# => x"fc",
        16#7a6# => x"c4",
        16#7a7# => x"fc",
        16#7a8# => x"c4",
        16#7a9# => x"fc",
        16#7aa# => x"c4",
        16#7ab# => x"fc",
        16#7ac# => x"c4",
        16#7ad# => x"fc",
        16#7ae# => x"c4",
        16#7af# => x"fc",
        16#7b0# => x"88",
        16#7b1# => x"f9",
        16#7b2# => x"88",
        16#7b3# => x"f9",
        16#7b4# => x"88",
        16#7b5# => x"f9",
        16#7b6# => x"36",
        16#7b7# => x"80",
        16#7b8# => x"ff",
        16#7b9# => x"4c",
        16#7ba# => x"c4",
        16#7bb# => x"fc",
        16#7bc# => x"4c",
        16#7bd# => x"c4",
        16#7be# => x"fc",
        16#7bf# => x"4c",
        16#7c0# => x"c4",
        16#7c1# => x"fc",
        16#7c2# => x"4c",
        16#7c3# => x"c4",
        16#7c4# => x"fc",
        16#7c5# => x"4c",
        16#7c6# => x"c4",
        16#7c7# => x"fc",
        16#7c8# => x"4c",
        16#7c9# => x"77",
        16#7ca# => x"f9",
        16#7cb# => x"4c",
        16#7cc# => x"6d",
        16#7cd# => x"f9",
        16#7ce# => x"6c",
        16#7cf# => x"1c",
        16#7d0# => x"02",
        16#7d1# => x"6c",
        16#7d2# => x"1a",
        16#7d3# => x"02",
        16#7d4# => x"6c",
        16#7d5# => x"18",
        16#7d6# => x"02",
        16#7d7# => x"6c",
        16#7d8# => x"16",
        16#7d9# => x"02",
        16#7da# => x"6c",
        16#7db# => x"14",
        16#7dc# => x"02",
        16#7dd# => x"6c",
        16#7de# => x"12",
        16#7df# => x"02",
        16#7e0# => x"6c",
        16#7e1# => x"10",
        16#7e2# => x"02",
        16#7e3# => x"c9",
        16#7e4# => x"0d",
        16#7e5# => x"d0",
        16#7e6# => x"07",
        16#7e7# => x"a9",
        16#7e8# => x"0a",
        16#7e9# => x"20",
        16#7ea# => x"ee",
        16#7eb# => x"ff",
        16#7ec# => x"a9",
        16#7ed# => x"0d",
        16#7ee# => x"6c",
        16#7ef# => x"0e",
        16#7f0# => x"02",
        16#7f1# => x"6c",
        16#7f2# => x"0c",
        16#7f3# => x"02",
        16#7f4# => x"6c",
        16#7f5# => x"0a",
        16#7f6# => x"02",
        16#7f7# => x"6c",
        16#7f8# => x"08",
        16#7f9# => x"02",
        16#7fa# => x"0d",
        16#7fb# => x"fe",
        16#7fc# => x"00",
        16#7fd# => x"f8",
        16#7fe# => x"f2",
        16#7ff# => x"fc"
        );

    attribute ram_style        : string;

    attribute ram_style of RAM : signal is "distributed";

begin

    process (CLK)
    begin
        if rising_edge(CLK) then
            DATA <= RAM(conv_integer(ADDR));            
        end if;
    end process;
    
end RTL;



