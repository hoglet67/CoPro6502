library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tuberom_65c102_banner is
    port (
        CLK  : in  std_logic;
        ADDR : in  std_logic_vector(10 downto 0);
        SW   : in  std_logic_vector(1 downto 0);
        DATA : out std_logic_vector(7 downto 0)
        );
end;

architecture RTL of tuberom_65c102_banner is

    signal rom_addr : std_logic_vector(11 downto 0);

    signal digit1 : std_logic_vector(7 downto 0);
    signal digit2 : std_logic_vector(7 downto 0);
    
begin

    p_addr : process(ADDR)
    begin
        rom_addr              <= (others => '0');
        rom_addr(10 downto 0) <= ADDR;
    end process;

    -- Original: Acorn TUBE 65C102 Co-Processor
    -- Updated:  Acorn TUBE 32Mhz 65C102 Co-Pro
    
    digit1 <= x"33" when SW = "00" else
              x"31" when SW = "01" else
              x"30"; 

    digit2 <= x"32" when SW = "00" else
              x"36" when SW = "01" else
              x"38" when SW = "10" else
              x"34";

    p_rom : process
    begin
        wait until rising_edge(CLK);
        DATA <= (others => '0');
        case rom_addr is
            when x"000" => DATA <= x"A2";
            when x"001" => DATA <= x"00";
            when x"002" => DATA <= x"BD";
            when x"003" => DATA <= x"00";
            when x"004" => DATA <= x"FF";
            when x"005" => DATA <= x"9D";
            when x"006" => DATA <= x"00";
            when x"007" => DATA <= x"FF";
            when x"008" => DATA <= x"CA";
            when x"009" => DATA <= x"D0";
            when x"00A" => DATA <= x"F7";
            when x"00B" => DATA <= x"A2";
            when x"00C" => DATA <= x"36";
            when x"00D" => DATA <= x"BD";
            when x"00E" => DATA <= x"80";
            when x"00F" => DATA <= x"FF";
            when x"010" => DATA <= x"9D";
            when x"011" => DATA <= x"00";
            when x"012" => DATA <= x"02";
            when x"013" => DATA <= x"CA";
            when x"014" => DATA <= x"10";
            when x"015" => DATA <= x"F7";
            when x"016" => DATA <= x"9A";
            when x"017" => DATA <= x"A2";
            when x"018" => DATA <= x"F0";
            when x"019" => DATA <= x"BD";
            when x"01A" => DATA <= x"FF";
            when x"01B" => DATA <= x"FD";
            when x"01C" => DATA <= x"9D";
            when x"01D" => DATA <= x"FF";
            when x"01E" => DATA <= x"FD";
            when x"01F" => DATA <= x"CA";
            when x"020" => DATA <= x"D0";
            when x"021" => DATA <= x"F7";
            when x"022" => DATA <= x"A0";
            when x"023" => DATA <= x"00";
            when x"024" => DATA <= x"84";
            when x"025" => DATA <= x"F8";
            when x"026" => DATA <= x"A9";
            when x"027" => DATA <= x"F8";
            when x"028" => DATA <= x"85";
            when x"029" => DATA <= x"F9";
            when x"02A" => DATA <= x"B1";
            when x"02B" => DATA <= x"F8";
            when x"02C" => DATA <= x"91";
            when x"02D" => DATA <= x"F8";
            when x"02E" => DATA <= x"C8";
            when x"02F" => DATA <= x"D0";
            when x"030" => DATA <= x"F9";
            when x"031" => DATA <= x"E6";
            when x"032" => DATA <= x"F9";
            when x"033" => DATA <= x"A5";
            when x"034" => DATA <= x"F9";
            when x"035" => DATA <= x"C9";
            when x"036" => DATA <= x"FE";
            when x"037" => DATA <= x"D0";
            when x"038" => DATA <= x"F1";
            when x"039" => DATA <= x"A2";
            when x"03A" => DATA <= x"10";
            when x"03B" => DATA <= x"BD";
            when x"03C" => DATA <= x"59";
            when x"03D" => DATA <= x"F8";
            when x"03E" => DATA <= x"9D";
            when x"03F" => DATA <= x"00";
            when x"040" => DATA <= x"01";
            when x"041" => DATA <= x"CA";
            when x"042" => DATA <= x"10";
            when x"043" => DATA <= x"F7";
            when x"044" => DATA <= x"A5";
            when x"045" => DATA <= x"EE";
            when x"046" => DATA <= x"85";
            when x"047" => DATA <= x"F6";
            when x"048" => DATA <= x"A5";
            when x"049" => DATA <= x"EF";
            when x"04A" => DATA <= x"85";
            when x"04B" => DATA <= x"F7";
            when x"04C" => DATA <= x"A9";
            when x"04D" => DATA <= x"00";
            when x"04E" => DATA <= x"85";
            when x"04F" => DATA <= x"FF";
            when x"050" => DATA <= x"85";
            when x"051" => DATA <= x"F2";
            when x"052" => DATA <= x"A9";
            when x"053" => DATA <= x"F8";
            when x"054" => DATA <= x"85";
            when x"055" => DATA <= x"F3";
            when x"056" => DATA <= x"4C";
            when x"057" => DATA <= x"00";
            when x"058" => DATA <= x"01";
            when x"059" => DATA <= x"AD";
            when x"05A" => DATA <= x"F8";
            when x"05B" => DATA <= x"FE";
            when x"05C" => DATA <= x"58";
            when x"05D" => DATA <= x"4C";
            when x"05E" => DATA <= x"60";
            when x"05F" => DATA <= x"F8";
            when x"060" => DATA <= x"20";
            when x"061" => DATA <= x"A5";
            when x"062" => DATA <= x"FE";
            when x"063" => DATA <= x"0A";
            when x"064" => DATA <= x"41";
            when x"065" => DATA <= x"63";
            when x"066" => DATA <= x"6F";
            when x"067" => DATA <= x"72";
            when x"068" => DATA <= x"6E";
            when x"069" => DATA <= x"20";
            when x"06A" => DATA <= x"54";
            when x"06B" => DATA <= x"55";
            when x"06C" => DATA <= x"42";
            when x"06D" => DATA <= x"45";
            when x"06E" => DATA <= x"20";
            when x"06F" => DATA <= digit1;
            when x"070" => DATA <= digit2;
            when x"071" => DATA <= x"4D";
            when x"072" => DATA <= x"68";
            when x"073" => DATA <= x"7A";
            when x"074" => DATA <= x"20";
            when x"075" => DATA <= x"36";
            when x"076" => DATA <= x"35";
            when x"077" => DATA <= x"43";
            when x"078" => DATA <= x"31";
            when x"079" => DATA <= x"30";
            when x"07A" => DATA <= x"32";
            when x"07B" => DATA <= x"20";
            when x"07C" => DATA <= x"43";
            when x"07D" => DATA <= x"6F";
            when x"07E" => DATA <= x"2D";
            when x"07F" => DATA <= x"50";
            when x"080" => DATA <= x"72";
            when x"081" => DATA <= x"6F";
            when x"082" => DATA <= x"0A";
            when x"083" => DATA <= x"0A";
            when x"084" => DATA <= x"0D";
            when x"085" => DATA <= x"00";
            when x"086" => DATA <= x"EA";
            when x"087" => DATA <= x"A9";
            when x"088" => DATA <= x"98";
            when x"089" => DATA <= x"8D";
            when x"08A" => DATA <= x"5E";
            when x"08B" => DATA <= x"F8";
            when x"08C" => DATA <= x"A9";
            when x"08D" => DATA <= x"F8";
            when x"08E" => DATA <= x"8D";
            when x"08F" => DATA <= x"5F";
            when x"090" => DATA <= x"F8";
            when x"091" => DATA <= x"20";
            when x"092" => DATA <= x"80";
            when x"093" => DATA <= x"F9";
            when x"094" => DATA <= x"C9";
            when x"095" => DATA <= x"80";
            when x"096" => DATA <= x"F0";
            when x"097" => DATA <= x"28";
            when x"098" => DATA <= x"A9";
            when x"099" => DATA <= x"2A";
            when x"09A" => DATA <= x"20";
            when x"09B" => DATA <= x"EE";
            when x"09C" => DATA <= x"FF";
            when x"09D" => DATA <= x"A2";
            when x"09E" => DATA <= x"68";
            when x"09F" => DATA <= x"A0";
            when x"0A0" => DATA <= x"F9";
            when x"0A1" => DATA <= x"A9";
            when x"0A2" => DATA <= x"00";
            when x"0A3" => DATA <= x"20";
            when x"0A4" => DATA <= x"F1";
            when x"0A5" => DATA <= x"FF";
            when x"0A6" => DATA <= x"B0";
            when x"0A7" => DATA <= x"0A";
            when x"0A8" => DATA <= x"A2";
            when x"0A9" => DATA <= x"36";
            when x"0AA" => DATA <= x"A0";
            when x"0AB" => DATA <= x"02";
            when x"0AC" => DATA <= x"20";
            when x"0AD" => DATA <= x"F7";
            when x"0AE" => DATA <= x"FF";
            when x"0AF" => DATA <= x"4C";
            when x"0B0" => DATA <= x"98";
            when x"0B1" => DATA <= x"F8";
            when x"0B2" => DATA <= x"A9";
            when x"0B3" => DATA <= x"7E";
            when x"0B4" => DATA <= x"20";
            when x"0B5" => DATA <= x"F4";
            when x"0B6" => DATA <= x"FF";
            when x"0B7" => DATA <= x"00";
            when x"0B8" => DATA <= x"11";
            when x"0B9" => DATA <= x"45";
            when x"0BA" => DATA <= x"73";
            when x"0BB" => DATA <= x"63";
            when x"0BC" => DATA <= x"61";
            when x"0BD" => DATA <= x"70";
            when x"0BE" => DATA <= x"65";
            when x"0BF" => DATA <= x"00";
            when x"0C0" => DATA <= x"A5";
            when x"0C1" => DATA <= x"F6";
            when x"0C2" => DATA <= x"85";
            when x"0C3" => DATA <= x"EE";
            when x"0C4" => DATA <= x"85";
            when x"0C5" => DATA <= x"F2";
            when x"0C6" => DATA <= x"A5";
            when x"0C7" => DATA <= x"F7";
            when x"0C8" => DATA <= x"85";
            when x"0C9" => DATA <= x"EF";
            when x"0CA" => DATA <= x"85";
            when x"0CB" => DATA <= x"F3";
            when x"0CC" => DATA <= x"A0";
            when x"0CD" => DATA <= x"07";
            when x"0CE" => DATA <= x"B1";
            when x"0CF" => DATA <= x"EE";
            when x"0D0" => DATA <= x"D8";
            when x"0D1" => DATA <= x"18";
            when x"0D2" => DATA <= x"65";
            when x"0D3" => DATA <= x"EE";
            when x"0D4" => DATA <= x"85";
            when x"0D5" => DATA <= x"FD";
            when x"0D6" => DATA <= x"A9";
            when x"0D7" => DATA <= x"00";
            when x"0D8" => DATA <= x"65";
            when x"0D9" => DATA <= x"EF";
            when x"0DA" => DATA <= x"85";
            when x"0DB" => DATA <= x"FE";
            when x"0DC" => DATA <= x"A0";
            when x"0DD" => DATA <= x"00";
            when x"0DE" => DATA <= x"B1";
            when x"0DF" => DATA <= x"FD";
            when x"0E0" => DATA <= x"D0";
            when x"0E1" => DATA <= x"23";
            when x"0E2" => DATA <= x"C8";
            when x"0E3" => DATA <= x"B1";
            when x"0E4" => DATA <= x"FD";
            when x"0E5" => DATA <= x"C9";
            when x"0E6" => DATA <= x"28";
            when x"0E7" => DATA <= x"D0";
            when x"0E8" => DATA <= x"1C";
            when x"0E9" => DATA <= x"C8";
            when x"0EA" => DATA <= x"B1";
            when x"0EB" => DATA <= x"FD";
            when x"0EC" => DATA <= x"C9";
            when x"0ED" => DATA <= x"43";
            when x"0EE" => DATA <= x"D0";
            when x"0EF" => DATA <= x"15";
            when x"0F0" => DATA <= x"C8";
            when x"0F1" => DATA <= x"B1";
            when x"0F2" => DATA <= x"FD";
            when x"0F3" => DATA <= x"C9";
            when x"0F4" => DATA <= x"29";
            when x"0F5" => DATA <= x"D0";
            when x"0F6" => DATA <= x"0E";
            when x"0F7" => DATA <= x"A0";
            when x"0F8" => DATA <= x"06";
            when x"0F9" => DATA <= x"B1";
            when x"0FA" => DATA <= x"EE";
            when x"0FB" => DATA <= x"29";
            when x"0FC" => DATA <= x"4F";
            when x"0FD" => DATA <= x"C9";
            when x"0FE" => DATA <= x"40";
            when x"0FF" => DATA <= x"90";
            when x"100" => DATA <= x"09";
            when x"101" => DATA <= x"29";
            when x"102" => DATA <= x"0D";
            when x"103" => DATA <= x"D0";
            when x"104" => DATA <= x"28";
            when x"105" => DATA <= x"A9";
            when x"106" => DATA <= x"01";
            when x"107" => DATA <= x"6C";
            when x"108" => DATA <= x"F2";
            when x"109" => DATA <= x"00";
            when x"10A" => DATA <= x"A9";
            when x"10B" => DATA <= x"50";
            when x"10C" => DATA <= x"8D";
            when x"10D" => DATA <= x"02";
            when x"10E" => DATA <= x"02";
            when x"10F" => DATA <= x"A9";
            when x"110" => DATA <= x"F9";
            when x"111" => DATA <= x"8D";
            when x"112" => DATA <= x"03";
            when x"113" => DATA <= x"02";
            when x"114" => DATA <= x"00";
            when x"115" => DATA <= x"00";
            when x"116" => DATA <= x"54";
            when x"117" => DATA <= x"68";
            when x"118" => DATA <= x"69";
            when x"119" => DATA <= x"73";
            when x"11A" => DATA <= x"20";
            when x"11B" => DATA <= x"69";
            when x"11C" => DATA <= x"73";
            when x"11D" => DATA <= x"20";
            when x"11E" => DATA <= x"6E";
            when x"11F" => DATA <= x"6F";
            when x"120" => DATA <= x"74";
            when x"121" => DATA <= x"20";
            when x"122" => DATA <= x"61";
            when x"123" => DATA <= x"20";
            when x"124" => DATA <= x"6C";
            when x"125" => DATA <= x"61";
            when x"126" => DATA <= x"6E";
            when x"127" => DATA <= x"67";
            when x"128" => DATA <= x"75";
            when x"129" => DATA <= x"61";
            when x"12A" => DATA <= x"67";
            when x"12B" => DATA <= x"65";
            when x"12C" => DATA <= x"00";
            when x"12D" => DATA <= x"A9";
            when x"12E" => DATA <= x"50";
            when x"12F" => DATA <= x"8D";
            when x"130" => DATA <= x"02";
            when x"131" => DATA <= x"02";
            when x"132" => DATA <= x"A9";
            when x"133" => DATA <= x"F9";
            when x"134" => DATA <= x"8D";
            when x"135" => DATA <= x"03";
            when x"136" => DATA <= x"02";
            when x"137" => DATA <= x"00";
            when x"138" => DATA <= x"00";
            when x"139" => DATA <= x"49";
            when x"13A" => DATA <= x"20";
            when x"13B" => DATA <= x"63";
            when x"13C" => DATA <= x"61";
            when x"13D" => DATA <= x"6E";
            when x"13E" => DATA <= x"6E";
            when x"13F" => DATA <= x"6F";
            when x"140" => DATA <= x"74";
            when x"141" => DATA <= x"20";
            when x"142" => DATA <= x"72";
            when x"143" => DATA <= x"75";
            when x"144" => DATA <= x"6E";
            when x"145" => DATA <= x"20";
            when x"146" => DATA <= x"74";
            when x"147" => DATA <= x"68";
            when x"148" => DATA <= x"69";
            when x"149" => DATA <= x"73";
            when x"14A" => DATA <= x"20";
            when x"14B" => DATA <= x"63";
            when x"14C" => DATA <= x"6F";
            when x"14D" => DATA <= x"64";
            when x"14E" => DATA <= x"65";
            when x"14F" => DATA <= x"00";
            when x"150" => DATA <= x"A2";
            when x"151" => DATA <= x"FF";
            when x"152" => DATA <= x"9A";
            when x"153" => DATA <= x"20";
            when x"154" => DATA <= x"E7";
            when x"155" => DATA <= x"FF";
            when x"156" => DATA <= x"A0";
            when x"157" => DATA <= x"01";
            when x"158" => DATA <= x"B1";
            when x"159" => DATA <= x"FD";
            when x"15A" => DATA <= x"F0";
            when x"15B" => DATA <= x"06";
            when x"15C" => DATA <= x"20";
            when x"15D" => DATA <= x"EE";
            when x"15E" => DATA <= x"FF";
            when x"15F" => DATA <= x"C8";
            when x"160" => DATA <= x"D0";
            when x"161" => DATA <= x"F6";
            when x"162" => DATA <= x"20";
            when x"163" => DATA <= x"E7";
            when x"164" => DATA <= x"FF";
            when x"165" => DATA <= x"4C";
            when x"166" => DATA <= x"98";
            when x"167" => DATA <= x"F8";
            when x"168" => DATA <= x"36";
            when x"169" => DATA <= x"02";
            when x"16A" => DATA <= x"CA";
            when x"16B" => DATA <= x"20";
            when x"16C" => DATA <= x"FF";
            when x"16D" => DATA <= x"2C";
            when x"16E" => DATA <= x"F8";
            when x"16F" => DATA <= x"FE";
            when x"170" => DATA <= x"EA";
            when x"171" => DATA <= x"50";
            when x"172" => DATA <= x"FA";
            when x"173" => DATA <= x"8D";
            when x"174" => DATA <= x"F9";
            when x"175" => DATA <= x"FE";
            when x"176" => DATA <= x"60";
            when x"177" => DATA <= x"A9";
            when x"178" => DATA <= x"00";
            when x"179" => DATA <= x"20";
            when x"17A" => DATA <= x"57";
            when x"17B" => DATA <= x"FC";
            when x"17C" => DATA <= x"20";
            when x"17D" => DATA <= x"80";
            when x"17E" => DATA <= x"F9";
            when x"17F" => DATA <= x"0A";
            when x"180" => DATA <= x"2C";
            when x"181" => DATA <= x"FA";
            when x"182" => DATA <= x"FE";
            when x"183" => DATA <= x"10";
            when x"184" => DATA <= x"FB";
            when x"185" => DATA <= x"AD";
            when x"186" => DATA <= x"FB";
            when x"187" => DATA <= x"FE";
            when x"188" => DATA <= x"60";
            when x"189" => DATA <= x"C8";
            when x"18A" => DATA <= x"B1";
            when x"18B" => DATA <= x"F8";
            when x"18C" => DATA <= x"C9";
            when x"18D" => DATA <= x"20";
            when x"18E" => DATA <= x"F0";
            when x"18F" => DATA <= x"F9";
            when x"190" => DATA <= x"60";
            when x"191" => DATA <= x"A2";
            when x"192" => DATA <= x"00";
            when x"193" => DATA <= x"86";
            when x"194" => DATA <= x"F0";
            when x"195" => DATA <= x"86";
            when x"196" => DATA <= x"F1";
            when x"197" => DATA <= x"B1";
            when x"198" => DATA <= x"F8";
            when x"199" => DATA <= x"C9";
            when x"19A" => DATA <= x"30";
            when x"19B" => DATA <= x"90";
            when x"19C" => DATA <= x"1F";
            when x"19D" => DATA <= x"C9";
            when x"19E" => DATA <= x"3A";
            when x"19F" => DATA <= x"90";
            when x"1A0" => DATA <= x"0A";
            when x"1A1" => DATA <= x"29";
            when x"1A2" => DATA <= x"DF";
            when x"1A3" => DATA <= x"E9";
            when x"1A4" => DATA <= x"07";
            when x"1A5" => DATA <= x"90";
            when x"1A6" => DATA <= x"15";
            when x"1A7" => DATA <= x"C9";
            when x"1A8" => DATA <= x"40";
            when x"1A9" => DATA <= x"B0";
            when x"1AA" => DATA <= x"11";
            when x"1AB" => DATA <= x"0A";
            when x"1AC" => DATA <= x"0A";
            when x"1AD" => DATA <= x"0A";
            when x"1AE" => DATA <= x"0A";
            when x"1AF" => DATA <= x"A2";
            when x"1B0" => DATA <= x"03";
            when x"1B1" => DATA <= x"0A";
            when x"1B2" => DATA <= x"26";
            when x"1B3" => DATA <= x"F0";
            when x"1B4" => DATA <= x"26";
            when x"1B5" => DATA <= x"F1";
            when x"1B6" => DATA <= x"CA";
            when x"1B7" => DATA <= x"10";
            when x"1B8" => DATA <= x"F8";
            when x"1B9" => DATA <= x"C8";
            when x"1BA" => DATA <= x"D0";
            when x"1BB" => DATA <= x"DB";
            when x"1BC" => DATA <= x"60";
            when x"1BD" => DATA <= x"86";
            when x"1BE" => DATA <= x"F8";
            when x"1BF" => DATA <= x"84";
            when x"1C0" => DATA <= x"F9";
            when x"1C1" => DATA <= x"A0";
            when x"1C2" => DATA <= x"00";
            when x"1C3" => DATA <= x"2C";
            when x"1C4" => DATA <= x"FA";
            when x"1C5" => DATA <= x"FE";
            when x"1C6" => DATA <= x"50";
            when x"1C7" => DATA <= x"FB";
            when x"1C8" => DATA <= x"B1";
            when x"1C9" => DATA <= x"F8";
            when x"1CA" => DATA <= x"8D";
            when x"1CB" => DATA <= x"FB";
            when x"1CC" => DATA <= x"FE";
            when x"1CD" => DATA <= x"C8";
            when x"1CE" => DATA <= x"C9";
            when x"1CF" => DATA <= x"0D";
            when x"1D0" => DATA <= x"D0";
            when x"1D1" => DATA <= x"F1";
            when x"1D2" => DATA <= x"A4";
            when x"1D3" => DATA <= x"F9";
            when x"1D4" => DATA <= x"60";
            when x"1D5" => DATA <= x"48";
            when x"1D6" => DATA <= x"86";
            when x"1D7" => DATA <= x"F8";
            when x"1D8" => DATA <= x"84";
            when x"1D9" => DATA <= x"F9";
            when x"1DA" => DATA <= x"A0";
            when x"1DB" => DATA <= x"00";
            when x"1DC" => DATA <= x"20";
            when x"1DD" => DATA <= x"8A";
            when x"1DE" => DATA <= x"F9";
            when x"1DF" => DATA <= x"C8";
            when x"1E0" => DATA <= x"C9";
            when x"1E1" => DATA <= x"2A";
            when x"1E2" => DATA <= x"F0";
            when x"1E3" => DATA <= x"F8";
            when x"1E4" => DATA <= x"29";
            when x"1E5" => DATA <= x"DF";
            when x"1E6" => DATA <= x"AA";
            when x"1E7" => DATA <= x"B1";
            when x"1E8" => DATA <= x"F8";
            when x"1E9" => DATA <= x"E0";
            when x"1EA" => DATA <= x"47";
            when x"1EB" => DATA <= x"F0";
            when x"1EC" => DATA <= x"5E";
            when x"1ED" => DATA <= x"E0";
            when x"1EE" => DATA <= x"48";
            when x"1EF" => DATA <= x"D0";
            when x"1F0" => DATA <= x"49";
            when x"1F1" => DATA <= x"C9";
            when x"1F2" => DATA <= x"2E";
            when x"1F3" => DATA <= x"F0";
            when x"1F4" => DATA <= x"2D";
            when x"1F5" => DATA <= x"29";
            when x"1F6" => DATA <= x"DF";
            when x"1F7" => DATA <= x"C9";
            when x"1F8" => DATA <= x"45";
            when x"1F9" => DATA <= x"D0";
            when x"1FA" => DATA <= x"3F";
            when x"1FB" => DATA <= x"C8";
            when x"1FC" => DATA <= x"B1";
            when x"1FD" => DATA <= x"F8";
            when x"1FE" => DATA <= x"C9";
            when x"1FF" => DATA <= x"2E";
            when x"200" => DATA <= x"F0";
            when x"201" => DATA <= x"20";
            when x"202" => DATA <= x"29";
            when x"203" => DATA <= x"DF";
            when x"204" => DATA <= x"C9";
            when x"205" => DATA <= x"4C";
            when x"206" => DATA <= x"D0";
            when x"207" => DATA <= x"32";
            when x"208" => DATA <= x"C8";
            when x"209" => DATA <= x"B1";
            when x"20A" => DATA <= x"F8";
            when x"20B" => DATA <= x"C9";
            when x"20C" => DATA <= x"2E";
            when x"20D" => DATA <= x"F0";
            when x"20E" => DATA <= x"13";
            when x"20F" => DATA <= x"29";
            when x"210" => DATA <= x"DF";
            when x"211" => DATA <= x"C9";
            when x"212" => DATA <= x"50";
            when x"213" => DATA <= x"D0";
            when x"214" => DATA <= x"25";
            when x"215" => DATA <= x"C8";
            when x"216" => DATA <= x"B1";
            when x"217" => DATA <= x"F8";
            when x"218" => DATA <= x"29";
            when x"219" => DATA <= x"DF";
            when x"21A" => DATA <= x"C9";
            when x"21B" => DATA <= x"41";
            when x"21C" => DATA <= x"90";
            when x"21D" => DATA <= x"04";
            when x"21E" => DATA <= x"C9";
            when x"21F" => DATA <= x"5B";
            when x"220" => DATA <= x"90";
            when x"221" => DATA <= x"18";
            when x"222" => DATA <= x"20";
            when x"223" => DATA <= x"A5";
            when x"224" => DATA <= x"FE";
            when x"225" => DATA <= x"0A";
            when x"226" => DATA <= x"0D";
            when x"227" => DATA <= x"36";
            when x"228" => DATA <= x"35";
            when x"229" => DATA <= x"43";
            when x"22A" => DATA <= x"31";
            when x"22B" => DATA <= x"30";
            when x"22C" => DATA <= x"32";
            when x"22D" => DATA <= x"20";
            when x"22E" => DATA <= x"54";
            when x"22F" => DATA <= x"55";
            when x"230" => DATA <= x"42";
            when x"231" => DATA <= x"45";
            when x"232" => DATA <= x"20";
            when x"233" => DATA <= x"31";
            when x"234" => DATA <= x"2E";
            when x"235" => DATA <= x"31";
            when x"236" => DATA <= x"30";
            when x"237" => DATA <= x"0A";
            when x"238" => DATA <= x"0D";
            when x"239" => DATA <= x"EA";
            when x"23A" => DATA <= x"A9";
            when x"23B" => DATA <= x"02";
            when x"23C" => DATA <= x"20";
            when x"23D" => DATA <= x"57";
            when x"23E" => DATA <= x"FC";
            when x"23F" => DATA <= x"20";
            when x"240" => DATA <= x"C1";
            when x"241" => DATA <= x"F9";
            when x"242" => DATA <= x"20";
            when x"243" => DATA <= x"80";
            when x"244" => DATA <= x"F9";
            when x"245" => DATA <= x"C9";
            when x"246" => DATA <= x"80";
            when x"247" => DATA <= x"F0";
            when x"248" => DATA <= x"20";
            when x"249" => DATA <= x"68";
            when x"24A" => DATA <= x"60";
            when x"24B" => DATA <= x"29";
            when x"24C" => DATA <= x"DF";
            when x"24D" => DATA <= x"C9";
            when x"24E" => DATA <= x"4F";
            when x"24F" => DATA <= x"D0";
            when x"250" => DATA <= x"E9";
            when x"251" => DATA <= x"20";
            when x"252" => DATA <= x"89";
            when x"253" => DATA <= x"F9";
            when x"254" => DATA <= x"20";
            when x"255" => DATA <= x"91";
            when x"256" => DATA <= x"F9";
            when x"257" => DATA <= x"20";
            when x"258" => DATA <= x"8A";
            when x"259" => DATA <= x"F9";
            when x"25A" => DATA <= x"C9";
            when x"25B" => DATA <= x"0D";
            when x"25C" => DATA <= x"D0";
            when x"25D" => DATA <= x"DC";
            when x"25E" => DATA <= x"8A";
            when x"25F" => DATA <= x"F0";
            when x"260" => DATA <= x"08";
            when x"261" => DATA <= x"A5";
            when x"262" => DATA <= x"F0";
            when x"263" => DATA <= x"85";
            when x"264" => DATA <= x"F6";
            when x"265" => DATA <= x"A5";
            when x"266" => DATA <= x"F1";
            when x"267" => DATA <= x"85";
            when x"268" => DATA <= x"F7";
            when x"269" => DATA <= x"A5";
            when x"26A" => DATA <= x"EF";
            when x"26B" => DATA <= x"48";
            when x"26C" => DATA <= x"A5";
            when x"26D" => DATA <= x"EE";
            when x"26E" => DATA <= x"48";
            when x"26F" => DATA <= x"20";
            when x"270" => DATA <= x"C0";
            when x"271" => DATA <= x"F8";
            when x"272" => DATA <= x"68";
            when x"273" => DATA <= x"85";
            when x"274" => DATA <= x"EE";
            when x"275" => DATA <= x"85";
            when x"276" => DATA <= x"F2";
            when x"277" => DATA <= x"68";
            when x"278" => DATA <= x"85";
            when x"279" => DATA <= x"EF";
            when x"27A" => DATA <= x"85";
            when x"27B" => DATA <= x"F3";
            when x"27C" => DATA <= x"68";
            when x"27D" => DATA <= x"60";
            when x"27E" => DATA <= x"F0";
            when x"27F" => DATA <= x"C2";
            when x"280" => DATA <= x"C9";
            when x"281" => DATA <= x"80";
            when x"282" => DATA <= x"B0";
            when x"283" => DATA <= x"25";
            when x"284" => DATA <= x"48";
            when x"285" => DATA <= x"A9";
            when x"286" => DATA <= x"04";
            when x"287" => DATA <= x"2C";
            when x"288" => DATA <= x"FA";
            when x"289" => DATA <= x"FE";
            when x"28A" => DATA <= x"50";
            when x"28B" => DATA <= x"FB";
            when x"28C" => DATA <= x"8D";
            when x"28D" => DATA <= x"FB";
            when x"28E" => DATA <= x"FE";
            when x"28F" => DATA <= x"2C";
            when x"290" => DATA <= x"FA";
            when x"291" => DATA <= x"FE";
            when x"292" => DATA <= x"50";
            when x"293" => DATA <= x"FB";
            when x"294" => DATA <= x"8E";
            when x"295" => DATA <= x"FB";
            when x"296" => DATA <= x"FE";
            when x"297" => DATA <= x"68";
            when x"298" => DATA <= x"2C";
            when x"299" => DATA <= x"FA";
            when x"29A" => DATA <= x"FE";
            when x"29B" => DATA <= x"50";
            when x"29C" => DATA <= x"FB";
            when x"29D" => DATA <= x"8D";
            when x"29E" => DATA <= x"FB";
            when x"29F" => DATA <= x"FE";
            when x"2A0" => DATA <= x"2C";
            when x"2A1" => DATA <= x"FA";
            when x"2A2" => DATA <= x"FE";
            when x"2A3" => DATA <= x"10";
            when x"2A4" => DATA <= x"FB";
            when x"2A5" => DATA <= x"AE";
            when x"2A6" => DATA <= x"FB";
            when x"2A7" => DATA <= x"FE";
            when x"2A8" => DATA <= x"60";
            when x"2A9" => DATA <= x"C9";
            when x"2AA" => DATA <= x"82";
            when x"2AB" => DATA <= x"F0";
            when x"2AC" => DATA <= x"5A";
            when x"2AD" => DATA <= x"C9";
            when x"2AE" => DATA <= x"83";
            when x"2AF" => DATA <= x"F0";
            when x"2B0" => DATA <= x"51";
            when x"2B1" => DATA <= x"C9";
            when x"2B2" => DATA <= x"84";
            when x"2B3" => DATA <= x"F0";
            when x"2B4" => DATA <= x"48";
            when x"2B5" => DATA <= x"48";
            when x"2B6" => DATA <= x"A9";
            when x"2B7" => DATA <= x"06";
            when x"2B8" => DATA <= x"2C";
            when x"2B9" => DATA <= x"FA";
            when x"2BA" => DATA <= x"FE";
            when x"2BB" => DATA <= x"50";
            when x"2BC" => DATA <= x"FB";
            when x"2BD" => DATA <= x"8D";
            when x"2BE" => DATA <= x"FB";
            when x"2BF" => DATA <= x"FE";
            when x"2C0" => DATA <= x"2C";
            when x"2C1" => DATA <= x"FA";
            when x"2C2" => DATA <= x"FE";
            when x"2C3" => DATA <= x"50";
            when x"2C4" => DATA <= x"FB";
            when x"2C5" => DATA <= x"8E";
            when x"2C6" => DATA <= x"FB";
            when x"2C7" => DATA <= x"FE";
            when x"2C8" => DATA <= x"2C";
            when x"2C9" => DATA <= x"FA";
            when x"2CA" => DATA <= x"FE";
            when x"2CB" => DATA <= x"50";
            when x"2CC" => DATA <= x"FB";
            when x"2CD" => DATA <= x"8C";
            when x"2CE" => DATA <= x"FB";
            when x"2CF" => DATA <= x"FE";
            when x"2D0" => DATA <= x"68";
            when x"2D1" => DATA <= x"2C";
            when x"2D2" => DATA <= x"FA";
            when x"2D3" => DATA <= x"FE";
            when x"2D4" => DATA <= x"50";
            when x"2D5" => DATA <= x"FB";
            when x"2D6" => DATA <= x"8D";
            when x"2D7" => DATA <= x"FB";
            when x"2D8" => DATA <= x"FE";
            when x"2D9" => DATA <= x"C9";
            when x"2DA" => DATA <= x"8E";
            when x"2DB" => DATA <= x"F0";
            when x"2DC" => DATA <= x"A1";
            when x"2DD" => DATA <= x"C9";
            when x"2DE" => DATA <= x"9D";
            when x"2DF" => DATA <= x"F0";
            when x"2E0" => DATA <= x"1B";
            when x"2E1" => DATA <= x"48";
            when x"2E2" => DATA <= x"2C";
            when x"2E3" => DATA <= x"FA";
            when x"2E4" => DATA <= x"FE";
            when x"2E5" => DATA <= x"10";
            when x"2E6" => DATA <= x"FB";
            when x"2E7" => DATA <= x"AD";
            when x"2E8" => DATA <= x"FB";
            when x"2E9" => DATA <= x"FE";
            when x"2EA" => DATA <= x"0A";
            when x"2EB" => DATA <= x"68";
            when x"2EC" => DATA <= x"2C";
            when x"2ED" => DATA <= x"FA";
            when x"2EE" => DATA <= x"FE";
            when x"2EF" => DATA <= x"10";
            when x"2F0" => DATA <= x"FB";
            when x"2F1" => DATA <= x"AC";
            when x"2F2" => DATA <= x"FB";
            when x"2F3" => DATA <= x"FE";
            when x"2F4" => DATA <= x"2C";
            when x"2F5" => DATA <= x"FA";
            when x"2F6" => DATA <= x"FE";
            when x"2F7" => DATA <= x"10";
            when x"2F8" => DATA <= x"FB";
            when x"2F9" => DATA <= x"AE";
            when x"2FA" => DATA <= x"FB";
            when x"2FB" => DATA <= x"FE";
            when x"2FC" => DATA <= x"60";
            when x"2FD" => DATA <= x"A6";
            when x"2FE" => DATA <= x"F2";
            when x"2FF" => DATA <= x"A4";
            when x"300" => DATA <= x"F3";
            when x"301" => DATA <= x"60";
            when x"302" => DATA <= x"A2";
            when x"303" => DATA <= x"00";
            when x"304" => DATA <= x"A0";
            when x"305" => DATA <= x"08";
            when x"306" => DATA <= x"60";
            when x"307" => DATA <= x"A2";
            when x"308" => DATA <= x"00";
            when x"309" => DATA <= x"A0";
            when x"30A" => DATA <= x"00";
            when x"30B" => DATA <= x"60";
            when x"30C" => DATA <= x"86";
            when x"30D" => DATA <= x"F8";
            when x"30E" => DATA <= x"84";
            when x"30F" => DATA <= x"F9";
            when x"310" => DATA <= x"A8";
            when x"311" => DATA <= x"F0";
            when x"312" => DATA <= x"71";
            when x"313" => DATA <= x"48";
            when x"314" => DATA <= x"A0";
            when x"315" => DATA <= x"08";
            when x"316" => DATA <= x"2C";
            when x"317" => DATA <= x"FA";
            when x"318" => DATA <= x"FE";
            when x"319" => DATA <= x"50";
            when x"31A" => DATA <= x"FB";
            when x"31B" => DATA <= x"8C";
            when x"31C" => DATA <= x"FB";
            when x"31D" => DATA <= x"FE";
            when x"31E" => DATA <= x"2C";
            when x"31F" => DATA <= x"FA";
            when x"320" => DATA <= x"FE";
            when x"321" => DATA <= x"50";
            when x"322" => DATA <= x"FB";
            when x"323" => DATA <= x"8D";
            when x"324" => DATA <= x"FB";
            when x"325" => DATA <= x"FE";
            when x"326" => DATA <= x"AA";
            when x"327" => DATA <= x"10";
            when x"328" => DATA <= x"08";
            when x"329" => DATA <= x"A0";
            when x"32A" => DATA <= x"00";
            when x"32B" => DATA <= x"B1";
            when x"32C" => DATA <= x"F8";
            when x"32D" => DATA <= x"A8";
            when x"32E" => DATA <= x"4C";
            when x"32F" => DATA <= x"3A";
            when x"330" => DATA <= x"FB";
            when x"331" => DATA <= x"BC";
            when x"332" => DATA <= x"C9";
            when x"333" => DATA <= x"FC";
            when x"334" => DATA <= x"E0";
            when x"335" => DATA <= x"15";
            when x"336" => DATA <= x"90";
            when x"337" => DATA <= x"02";
            when x"338" => DATA <= x"A0";
            when x"339" => DATA <= x"10";
            when x"33A" => DATA <= x"2C";
            when x"33B" => DATA <= x"FA";
            when x"33C" => DATA <= x"FE";
            when x"33D" => DATA <= x"50";
            when x"33E" => DATA <= x"FB";
            when x"33F" => DATA <= x"8C";
            when x"340" => DATA <= x"FB";
            when x"341" => DATA <= x"FE";
            when x"342" => DATA <= x"88";
            when x"343" => DATA <= x"30";
            when x"344" => DATA <= x"0D";
            when x"345" => DATA <= x"2C";
            when x"346" => DATA <= x"FA";
            when x"347" => DATA <= x"FE";
            when x"348" => DATA <= x"50";
            when x"349" => DATA <= x"FB";
            when x"34A" => DATA <= x"B1";
            when x"34B" => DATA <= x"F8";
            when x"34C" => DATA <= x"8D";
            when x"34D" => DATA <= x"FB";
            when x"34E" => DATA <= x"FE";
            when x"34F" => DATA <= x"88";
            when x"350" => DATA <= x"10";
            when x"351" => DATA <= x"F3";
            when x"352" => DATA <= x"8A";
            when x"353" => DATA <= x"10";
            when x"354" => DATA <= x"08";
            when x"355" => DATA <= x"A0";
            when x"356" => DATA <= x"01";
            when x"357" => DATA <= x"B1";
            when x"358" => DATA <= x"F8";
            when x"359" => DATA <= x"A8";
            when x"35A" => DATA <= x"4C";
            when x"35B" => DATA <= x"66";
            when x"35C" => DATA <= x"FB";
            when x"35D" => DATA <= x"BC";
            when x"35E" => DATA <= x"DD";
            when x"35F" => DATA <= x"FC";
            when x"360" => DATA <= x"E0";
            when x"361" => DATA <= x"15";
            when x"362" => DATA <= x"90";
            when x"363" => DATA <= x"02";
            when x"364" => DATA <= x"A0";
            when x"365" => DATA <= x"10";
            when x"366" => DATA <= x"2C";
            when x"367" => DATA <= x"FA";
            when x"368" => DATA <= x"FE";
            when x"369" => DATA <= x"50";
            when x"36A" => DATA <= x"FB";
            when x"36B" => DATA <= x"8C";
            when x"36C" => DATA <= x"FB";
            when x"36D" => DATA <= x"FE";
            when x"36E" => DATA <= x"88";
            when x"36F" => DATA <= x"30";
            when x"370" => DATA <= x"0D";
            when x"371" => DATA <= x"2C";
            when x"372" => DATA <= x"FA";
            when x"373" => DATA <= x"FE";
            when x"374" => DATA <= x"10";
            when x"375" => DATA <= x"FB";
            when x"376" => DATA <= x"AD";
            when x"377" => DATA <= x"FB";
            when x"378" => DATA <= x"FE";
            when x"379" => DATA <= x"91";
            when x"37A" => DATA <= x"F8";
            when x"37B" => DATA <= x"88";
            when x"37C" => DATA <= x"10";
            when x"37D" => DATA <= x"F3";
            when x"37E" => DATA <= x"A4";
            when x"37F" => DATA <= x"F9";
            when x"380" => DATA <= x"A6";
            when x"381" => DATA <= x"F8";
            when x"382" => DATA <= x"68";
            when x"383" => DATA <= x"60";
            when x"384" => DATA <= x"A9";
            when x"385" => DATA <= x"0A";
            when x"386" => DATA <= x"20";
            when x"387" => DATA <= x"57";
            when x"388" => DATA <= x"FC";
            when x"389" => DATA <= x"A0";
            when x"38A" => DATA <= x"04";
            when x"38B" => DATA <= x"2C";
            when x"38C" => DATA <= x"FA";
            when x"38D" => DATA <= x"FE";
            when x"38E" => DATA <= x"50";
            when x"38F" => DATA <= x"FB";
            when x"390" => DATA <= x"B1";
            when x"391" => DATA <= x"F8";
            when x"392" => DATA <= x"8D";
            when x"393" => DATA <= x"FB";
            when x"394" => DATA <= x"FE";
            when x"395" => DATA <= x"88";
            when x"396" => DATA <= x"C0";
            when x"397" => DATA <= x"01";
            when x"398" => DATA <= x"D0";
            when x"399" => DATA <= x"F1";
            when x"39A" => DATA <= x"A9";
            when x"39B" => DATA <= x"07";
            when x"39C" => DATA <= x"20";
            when x"39D" => DATA <= x"57";
            when x"39E" => DATA <= x"FC";
            when x"39F" => DATA <= x"B1";
            when x"3A0" => DATA <= x"F8";
            when x"3A1" => DATA <= x"48";
            when x"3A2" => DATA <= x"88";
            when x"3A3" => DATA <= x"2C";
            when x"3A4" => DATA <= x"FA";
            when x"3A5" => DATA <= x"FE";
            when x"3A6" => DATA <= x"50";
            when x"3A7" => DATA <= x"FB";
            when x"3A8" => DATA <= x"8C";
            when x"3A9" => DATA <= x"FB";
            when x"3AA" => DATA <= x"FE";
            when x"3AB" => DATA <= x"B1";
            when x"3AC" => DATA <= x"F8";
            when x"3AD" => DATA <= x"48";
            when x"3AE" => DATA <= x"A2";
            when x"3AF" => DATA <= x"FF";
            when x"3B0" => DATA <= x"20";
            when x"3B1" => DATA <= x"80";
            when x"3B2" => DATA <= x"F9";
            when x"3B3" => DATA <= x"C9";
            when x"3B4" => DATA <= x"80";
            when x"3B5" => DATA <= x"B0";
            when x"3B6" => DATA <= x"1D";
            when x"3B7" => DATA <= x"68";
            when x"3B8" => DATA <= x"85";
            when x"3B9" => DATA <= x"F8";
            when x"3BA" => DATA <= x"68";
            when x"3BB" => DATA <= x"85";
            when x"3BC" => DATA <= x"F9";
            when x"3BD" => DATA <= x"A0";
            when x"3BE" => DATA <= x"00";
            when x"3BF" => DATA <= x"2C";
            when x"3C0" => DATA <= x"FA";
            when x"3C1" => DATA <= x"FE";
            when x"3C2" => DATA <= x"10";
            when x"3C3" => DATA <= x"FB";
            when x"3C4" => DATA <= x"AD";
            when x"3C5" => DATA <= x"FB";
            when x"3C6" => DATA <= x"FE";
            when x"3C7" => DATA <= x"91";
            when x"3C8" => DATA <= x"F8";
            when x"3C9" => DATA <= x"C8";
            when x"3CA" => DATA <= x"C9";
            when x"3CB" => DATA <= x"0D";
            when x"3CC" => DATA <= x"D0";
            when x"3CD" => DATA <= x"F1";
            when x"3CE" => DATA <= x"A9";
            when x"3CF" => DATA <= x"00";
            when x"3D0" => DATA <= x"88";
            when x"3D1" => DATA <= x"18";
            when x"3D2" => DATA <= x"E8";
            when x"3D3" => DATA <= x"60";
            when x"3D4" => DATA <= x"68";
            when x"3D5" => DATA <= x"68";
            when x"3D6" => DATA <= x"A9";
            when x"3D7" => DATA <= x"00";
            when x"3D8" => DATA <= x"60";
            when x"3D9" => DATA <= x"48";
            when x"3DA" => DATA <= x"A9";
            when x"3DB" => DATA <= x"0C";
            when x"3DC" => DATA <= x"20";
            when x"3DD" => DATA <= x"57";
            when x"3DE" => DATA <= x"FC";
            when x"3DF" => DATA <= x"2C";
            when x"3E0" => DATA <= x"FA";
            when x"3E1" => DATA <= x"FE";
            when x"3E2" => DATA <= x"50";
            when x"3E3" => DATA <= x"FB";
            when x"3E4" => DATA <= x"8C";
            when x"3E5" => DATA <= x"FB";
            when x"3E6" => DATA <= x"FE";
            when x"3E7" => DATA <= x"B5";
            when x"3E8" => DATA <= x"03";
            when x"3E9" => DATA <= x"20";
            when x"3EA" => DATA <= x"57";
            when x"3EB" => DATA <= x"FC";
            when x"3EC" => DATA <= x"B5";
            when x"3ED" => DATA <= x"02";
            when x"3EE" => DATA <= x"20";
            when x"3EF" => DATA <= x"57";
            when x"3F0" => DATA <= x"FC";
            when x"3F1" => DATA <= x"B5";
            when x"3F2" => DATA <= x"01";
            when x"3F3" => DATA <= x"20";
            when x"3F4" => DATA <= x"57";
            when x"3F5" => DATA <= x"FC";
            when x"3F6" => DATA <= x"B5";
            when x"3F7" => DATA <= x"00";
            when x"3F8" => DATA <= x"20";
            when x"3F9" => DATA <= x"57";
            when x"3FA" => DATA <= x"FC";
            when x"3FB" => DATA <= x"68";
            when x"3FC" => DATA <= x"20";
            when x"3FD" => DATA <= x"57";
            when x"3FE" => DATA <= x"FC";
            when x"3FF" => DATA <= x"20";
            when x"400" => DATA <= x"80";
            when x"401" => DATA <= x"F9";
            when x"402" => DATA <= x"48";
            when x"403" => DATA <= x"20";
            when x"404" => DATA <= x"80";
            when x"405" => DATA <= x"F9";
            when x"406" => DATA <= x"95";
            when x"407" => DATA <= x"03";
            when x"408" => DATA <= x"20";
            when x"409" => DATA <= x"80";
            when x"40A" => DATA <= x"F9";
            when x"40B" => DATA <= x"95";
            when x"40C" => DATA <= x"02";
            when x"40D" => DATA <= x"20";
            when x"40E" => DATA <= x"80";
            when x"40F" => DATA <= x"F9";
            when x"410" => DATA <= x"95";
            when x"411" => DATA <= x"01";
            when x"412" => DATA <= x"20";
            when x"413" => DATA <= x"80";
            when x"414" => DATA <= x"F9";
            when x"415" => DATA <= x"95";
            when x"416" => DATA <= x"00";
            when x"417" => DATA <= x"68";
            when x"418" => DATA <= x"60";
            when x"419" => DATA <= x"48";
            when x"41A" => DATA <= x"A9";
            when x"41B" => DATA <= x"12";
            when x"41C" => DATA <= x"20";
            when x"41D" => DATA <= x"57";
            when x"41E" => DATA <= x"FC";
            when x"41F" => DATA <= x"68";
            when x"420" => DATA <= x"20";
            when x"421" => DATA <= x"57";
            when x"422" => DATA <= x"FC";
            when x"423" => DATA <= x"C9";
            when x"424" => DATA <= x"00";
            when x"425" => DATA <= x"D0";
            when x"426" => DATA <= x"0A";
            when x"427" => DATA <= x"48";
            when x"428" => DATA <= x"98";
            when x"429" => DATA <= x"20";
            when x"42A" => DATA <= x"57";
            when x"42B" => DATA <= x"FC";
            when x"42C" => DATA <= x"20";
            when x"42D" => DATA <= x"80";
            when x"42E" => DATA <= x"F9";
            when x"42F" => DATA <= x"68";
            when x"430" => DATA <= x"60";
            when x"431" => DATA <= x"20";
            when x"432" => DATA <= x"BD";
            when x"433" => DATA <= x"F9";
            when x"434" => DATA <= x"4C";
            when x"435" => DATA <= x"80";
            when x"436" => DATA <= x"F9";
            when x"437" => DATA <= x"A9";
            when x"438" => DATA <= x"0E";
            when x"439" => DATA <= x"20";
            when x"43A" => DATA <= x"57";
            when x"43B" => DATA <= x"FC";
            when x"43C" => DATA <= x"98";
            when x"43D" => DATA <= x"20";
            when x"43E" => DATA <= x"57";
            when x"43F" => DATA <= x"FC";
            when x"440" => DATA <= x"4C";
            when x"441" => DATA <= x"7C";
            when x"442" => DATA <= x"F9";
            when x"443" => DATA <= x"48";
            when x"444" => DATA <= x"A9";
            when x"445" => DATA <= x"10";
            when x"446" => DATA <= x"20";
            when x"447" => DATA <= x"57";
            when x"448" => DATA <= x"FC";
            when x"449" => DATA <= x"98";
            when x"44A" => DATA <= x"20";
            when x"44B" => DATA <= x"57";
            when x"44C" => DATA <= x"FC";
            when x"44D" => DATA <= x"68";
            when x"44E" => DATA <= x"20";
            when x"44F" => DATA <= x"57";
            when x"450" => DATA <= x"FC";
            when x"451" => DATA <= x"48";
            when x"452" => DATA <= x"20";
            when x"453" => DATA <= x"80";
            when x"454" => DATA <= x"F9";
            when x"455" => DATA <= x"68";
            when x"456" => DATA <= x"60";
            when x"457" => DATA <= x"2C";
            when x"458" => DATA <= x"FA";
            when x"459" => DATA <= x"FE";
            when x"45A" => DATA <= x"50";
            when x"45B" => DATA <= x"FB";
            when x"45C" => DATA <= x"8D";
            when x"45D" => DATA <= x"FB";
            when x"45E" => DATA <= x"FE";
            when x"45F" => DATA <= x"60";
            when x"460" => DATA <= x"84";
            when x"461" => DATA <= x"FB";
            when x"462" => DATA <= x"86";
            when x"463" => DATA <= x"FA";
            when x"464" => DATA <= x"48";
            when x"465" => DATA <= x"A9";
            when x"466" => DATA <= x"14";
            when x"467" => DATA <= x"20";
            when x"468" => DATA <= x"57";
            when x"469" => DATA <= x"FC";
            when x"46A" => DATA <= x"A0";
            when x"46B" => DATA <= x"11";
            when x"46C" => DATA <= x"B1";
            when x"46D" => DATA <= x"FA";
            when x"46E" => DATA <= x"20";
            when x"46F" => DATA <= x"57";
            when x"470" => DATA <= x"FC";
            when x"471" => DATA <= x"88";
            when x"472" => DATA <= x"C0";
            when x"473" => DATA <= x"01";
            when x"474" => DATA <= x"D0";
            when x"475" => DATA <= x"F6";
            when x"476" => DATA <= x"88";
            when x"477" => DATA <= x"B1";
            when x"478" => DATA <= x"FA";
            when x"479" => DATA <= x"AA";
            when x"47A" => DATA <= x"C8";
            when x"47B" => DATA <= x"B1";
            when x"47C" => DATA <= x"FA";
            when x"47D" => DATA <= x"A8";
            when x"47E" => DATA <= x"20";
            when x"47F" => DATA <= x"BD";
            when x"480" => DATA <= x"F9";
            when x"481" => DATA <= x"68";
            when x"482" => DATA <= x"20";
            when x"483" => DATA <= x"57";
            when x"484" => DATA <= x"FC";
            when x"485" => DATA <= x"20";
            when x"486" => DATA <= x"80";
            when x"487" => DATA <= x"F9";
            when x"488" => DATA <= x"48";
            when x"489" => DATA <= x"A0";
            when x"48A" => DATA <= x"11";
            when x"48B" => DATA <= x"20";
            when x"48C" => DATA <= x"80";
            when x"48D" => DATA <= x"F9";
            when x"48E" => DATA <= x"91";
            when x"48F" => DATA <= x"FA";
            when x"490" => DATA <= x"88";
            when x"491" => DATA <= x"C0";
            when x"492" => DATA <= x"01";
            when x"493" => DATA <= x"D0";
            when x"494" => DATA <= x"F6";
            when x"495" => DATA <= x"A4";
            when x"496" => DATA <= x"FB";
            when x"497" => DATA <= x"A6";
            when x"498" => DATA <= x"FA";
            when x"499" => DATA <= x"68";
            when x"49A" => DATA <= x"60";
            when x"49B" => DATA <= x"84";
            when x"49C" => DATA <= x"FB";
            when x"49D" => DATA <= x"86";
            when x"49E" => DATA <= x"FA";
            when x"49F" => DATA <= x"48";
            when x"4A0" => DATA <= x"A9";
            when x"4A1" => DATA <= x"16";
            when x"4A2" => DATA <= x"20";
            when x"4A3" => DATA <= x"57";
            when x"4A4" => DATA <= x"FC";
            when x"4A5" => DATA <= x"A0";
            when x"4A6" => DATA <= x"0C";
            when x"4A7" => DATA <= x"B1";
            when x"4A8" => DATA <= x"FA";
            when x"4A9" => DATA <= x"20";
            when x"4AA" => DATA <= x"57";
            when x"4AB" => DATA <= x"FC";
            when x"4AC" => DATA <= x"88";
            when x"4AD" => DATA <= x"10";
            when x"4AE" => DATA <= x"F8";
            when x"4AF" => DATA <= x"68";
            when x"4B0" => DATA <= x"20";
            when x"4B1" => DATA <= x"57";
            when x"4B2" => DATA <= x"FC";
            when x"4B3" => DATA <= x"A0";
            when x"4B4" => DATA <= x"0C";
            when x"4B5" => DATA <= x"20";
            when x"4B6" => DATA <= x"80";
            when x"4B7" => DATA <= x"F9";
            when x"4B8" => DATA <= x"91";
            when x"4B9" => DATA <= x"FA";
            when x"4BA" => DATA <= x"88";
            when x"4BB" => DATA <= x"10";
            when x"4BC" => DATA <= x"F8";
            when x"4BD" => DATA <= x"A4";
            when x"4BE" => DATA <= x"FB";
            when x"4BF" => DATA <= x"A6";
            when x"4C0" => DATA <= x"FA";
            when x"4C1" => DATA <= x"4C";
            when x"4C2" => DATA <= x"7C";
            when x"4C3" => DATA <= x"F9";
            when x"4C4" => DATA <= x"00";
            when x"4C5" => DATA <= x"FF";
            when x"4C6" => DATA <= x"42";
            when x"4C7" => DATA <= x"61";
            when x"4C8" => DATA <= x"64";
            when x"4C9" => DATA <= x"00";
            when x"4CA" => DATA <= x"00";
            when x"4CB" => DATA <= x"05";
            when x"4CC" => DATA <= x"00";
            when x"4CD" => DATA <= x"05";
            when x"4CE" => DATA <= x"04";
            when x"4CF" => DATA <= x"05";
            when x"4D0" => DATA <= x"08";
            when x"4D1" => DATA <= x"0E";
            when x"4D2" => DATA <= x"04";
            when x"4D3" => DATA <= x"01";
            when x"4D4" => DATA <= x"01";
            when x"4D5" => DATA <= x"05";
            when x"4D6" => DATA <= x"00";
            when x"4D7" => DATA <= x"01";
            when x"4D8" => DATA <= x"20";
            when x"4D9" => DATA <= x"10";
            when x"4DA" => DATA <= x"0D";
            when x"4DB" => DATA <= x"00";
            when x"4DC" => DATA <= x"04";
            when x"4DD" => DATA <= x"80";
            when x"4DE" => DATA <= x"05";
            when x"4DF" => DATA <= x"00";
            when x"4E0" => DATA <= x"05";
            when x"4E1" => DATA <= x"00";
            when x"4E2" => DATA <= x"05";
            when x"4E3" => DATA <= x"00";
            when x"4E4" => DATA <= x"00";
            when x"4E5" => DATA <= x"00";
            when x"4E6" => DATA <= x"05";
            when x"4E7" => DATA <= x"09";
            when x"4E8" => DATA <= x"05";
            when x"4E9" => DATA <= x"00";
            when x"4EA" => DATA <= x"08";
            when x"4EB" => DATA <= x"18";
            when x"4EC" => DATA <= x"00";
            when x"4ED" => DATA <= x"01";
            when x"4EE" => DATA <= x"0D";
            when x"4EF" => DATA <= x"80";
            when x"4F0" => DATA <= x"04";
            when x"4F1" => DATA <= x"80";
            when x"4F2" => DATA <= x"85";
            when x"4F3" => DATA <= x"FC";
            when x"4F4" => DATA <= x"68";
            when x"4F5" => DATA <= x"48";
            when x"4F6" => DATA <= x"29";
            when x"4F7" => DATA <= x"10";
            when x"4F8" => DATA <= x"D0";
            when x"4F9" => DATA <= x"10";
            when x"4FA" => DATA <= x"6C";
            when x"4FB" => DATA <= x"04";
            when x"4FC" => DATA <= x"02";
            when x"4FD" => DATA <= x"2C";
            when x"4FE" => DATA <= x"FE";
            when x"4FF" => DATA <= x"FE";
            when x"500" => DATA <= x"30";
            when x"501" => DATA <= x"4A";
            when x"502" => DATA <= x"2C";
            when x"503" => DATA <= x"F8";
            when x"504" => DATA <= x"FE";
            when x"505" => DATA <= x"30";
            when x"506" => DATA <= x"1E";
            when x"507" => DATA <= x"6C";
            when x"508" => DATA <= x"06";
            when x"509" => DATA <= x"02";
            when x"50A" => DATA <= x"8A";
            when x"50B" => DATA <= x"48";
            when x"50C" => DATA <= x"BA";
            when x"50D" => DATA <= x"BD";
            when x"50E" => DATA <= x"03";
            when x"50F" => DATA <= x"01";
            when x"510" => DATA <= x"D8";
            when x"511" => DATA <= x"38";
            when x"512" => DATA <= x"E9";
            when x"513" => DATA <= x"01";
            when x"514" => DATA <= x"85";
            when x"515" => DATA <= x"FD";
            when x"516" => DATA <= x"BD";
            when x"517" => DATA <= x"04";
            when x"518" => DATA <= x"01";
            when x"519" => DATA <= x"E9";
            when x"51A" => DATA <= x"00";
            when x"51B" => DATA <= x"85";
            when x"51C" => DATA <= x"FE";
            when x"51D" => DATA <= x"68";
            when x"51E" => DATA <= x"AA";
            when x"51F" => DATA <= x"A5";
            when x"520" => DATA <= x"FC";
            when x"521" => DATA <= x"58";
            when x"522" => DATA <= x"6C";
            when x"523" => DATA <= x"02";
            when x"524" => DATA <= x"02";
            when x"525" => DATA <= x"AD";
            when x"526" => DATA <= x"F9";
            when x"527" => DATA <= x"FE";
            when x"528" => DATA <= x"30";
            when x"529" => DATA <= x"1C";
            when x"52A" => DATA <= x"98";
            when x"52B" => DATA <= x"48";
            when x"52C" => DATA <= x"8A";
            when x"52D" => DATA <= x"48";
            when x"52E" => DATA <= x"20";
            when x"52F" => DATA <= x"8D";
            when x"530" => DATA <= x"FE";
            when x"531" => DATA <= x"A8";
            when x"532" => DATA <= x"20";
            when x"533" => DATA <= x"8D";
            when x"534" => DATA <= x"FE";
            when x"535" => DATA <= x"AA";
            when x"536" => DATA <= x"20";
            when x"537" => DATA <= x"8D";
            when x"538" => DATA <= x"FE";
            when x"539" => DATA <= x"20";
            when x"53A" => DATA <= x"43";
            when x"53B" => DATA <= x"FD";
            when x"53C" => DATA <= x"68";
            when x"53D" => DATA <= x"AA";
            when x"53E" => DATA <= x"68";
            when x"53F" => DATA <= x"A8";
            when x"540" => DATA <= x"A5";
            when x"541" => DATA <= x"FC";
            when x"542" => DATA <= x"40";
            when x"543" => DATA <= x"6C";
            when x"544" => DATA <= x"20";
            when x"545" => DATA <= x"02";
            when x"546" => DATA <= x"0A";
            when x"547" => DATA <= x"85";
            when x"548" => DATA <= x"FF";
            when x"549" => DATA <= x"A5";
            when x"54A" => DATA <= x"FC";
            when x"54B" => DATA <= x"40";
            when x"54C" => DATA <= x"AD";
            when x"54D" => DATA <= x"FF";
            when x"54E" => DATA <= x"FE";
            when x"54F" => DATA <= x"10";
            when x"550" => DATA <= x"21";
            when x"551" => DATA <= x"58";
            when x"552" => DATA <= x"2C";
            when x"553" => DATA <= x"FA";
            when x"554" => DATA <= x"FE";
            when x"555" => DATA <= x"10";
            when x"556" => DATA <= x"FB";
            when x"557" => DATA <= x"AD";
            when x"558" => DATA <= x"FB";
            when x"559" => DATA <= x"FE";
            when x"55A" => DATA <= x"A9";
            when x"55B" => DATA <= x"00";
            when x"55C" => DATA <= x"8D";
            when x"55D" => DATA <= x"36";
            when x"55E" => DATA <= x"02";
            when x"55F" => DATA <= x"A8";
            when x"560" => DATA <= x"20";
            when x"561" => DATA <= x"80";
            when x"562" => DATA <= x"F9";
            when x"563" => DATA <= x"8D";
            when x"564" => DATA <= x"37";
            when x"565" => DATA <= x"02";
            when x"566" => DATA <= x"C8";
            when x"567" => DATA <= x"20";
            when x"568" => DATA <= x"80";
            when x"569" => DATA <= x"F9";
            when x"56A" => DATA <= x"99";
            when x"56B" => DATA <= x"37";
            when x"56C" => DATA <= x"02";
            when x"56D" => DATA <= x"D0";
            when x"56E" => DATA <= x"F7";
            when x"56F" => DATA <= x"4C";
            when x"570" => DATA <= x"36";
            when x"571" => DATA <= x"02";
            when x"572" => DATA <= x"8D";
            when x"573" => DATA <= x"FA";
            when x"574" => DATA <= x"FF";
            when x"575" => DATA <= x"98";
            when x"576" => DATA <= x"48";
            when x"577" => DATA <= x"AC";
            when x"578" => DATA <= x"FA";
            when x"579" => DATA <= x"FF";
            when x"57A" => DATA <= x"B9";
            when x"57B" => DATA <= x"7D";
            when x"57C" => DATA <= x"FE";
            when x"57D" => DATA <= x"8D";
            when x"57E" => DATA <= x"FA";
            when x"57F" => DATA <= x"FF";
            when x"580" => DATA <= x"B9";
            when x"581" => DATA <= x"85";
            when x"582" => DATA <= x"FE";
            when x"583" => DATA <= x"8D";
            when x"584" => DATA <= x"FB";
            when x"585" => DATA <= x"FF";
            when x"586" => DATA <= x"B9";
            when x"587" => DATA <= x"6D";
            when x"588" => DATA <= x"FE";
            when x"589" => DATA <= x"85";
            when x"58A" => DATA <= x"F4";
            when x"58B" => DATA <= x"B9";
            when x"58C" => DATA <= x"75";
            when x"58D" => DATA <= x"FE";
            when x"58E" => DATA <= x"85";
            when x"58F" => DATA <= x"F5";
            when x"590" => DATA <= x"2C";
            when x"591" => DATA <= x"FE";
            when x"592" => DATA <= x"FE";
            when x"593" => DATA <= x"10";
            when x"594" => DATA <= x"FB";
            when x"595" => DATA <= x"AD";
            when x"596" => DATA <= x"FF";
            when x"597" => DATA <= x"FE";
            when x"598" => DATA <= x"C0";
            when x"599" => DATA <= x"05";
            when x"59A" => DATA <= x"F0";
            when x"59B" => DATA <= x"58";
            when x"59C" => DATA <= x"98";
            when x"59D" => DATA <= x"48";
            when x"59E" => DATA <= x"A0";
            when x"59F" => DATA <= x"01";
            when x"5A0" => DATA <= x"2C";
            when x"5A1" => DATA <= x"FE";
            when x"5A2" => DATA <= x"FE";
            when x"5A3" => DATA <= x"10";
            when x"5A4" => DATA <= x"FB";
            when x"5A5" => DATA <= x"AD";
            when x"5A6" => DATA <= x"FF";
            when x"5A7" => DATA <= x"FE";
            when x"5A8" => DATA <= x"2C";
            when x"5A9" => DATA <= x"FE";
            when x"5AA" => DATA <= x"FE";
            when x"5AB" => DATA <= x"10";
            when x"5AC" => DATA <= x"FB";
            when x"5AD" => DATA <= x"AD";
            when x"5AE" => DATA <= x"FF";
            when x"5AF" => DATA <= x"FE";
            when x"5B0" => DATA <= x"2C";
            when x"5B1" => DATA <= x"FE";
            when x"5B2" => DATA <= x"FE";
            when x"5B3" => DATA <= x"10";
            when x"5B4" => DATA <= x"FB";
            when x"5B5" => DATA <= x"AD";
            when x"5B6" => DATA <= x"FF";
            when x"5B7" => DATA <= x"FE";
            when x"5B8" => DATA <= x"91";
            when x"5B9" => DATA <= x"F4";
            when x"5BA" => DATA <= x"88";
            when x"5BB" => DATA <= x"2C";
            when x"5BC" => DATA <= x"FE";
            when x"5BD" => DATA <= x"FE";
            when x"5BE" => DATA <= x"10";
            when x"5BF" => DATA <= x"FB";
            when x"5C0" => DATA <= x"AD";
            when x"5C1" => DATA <= x"FF";
            when x"5C2" => DATA <= x"FE";
            when x"5C3" => DATA <= x"91";
            when x"5C4" => DATA <= x"F4";
            when x"5C5" => DATA <= x"2C";
            when x"5C6" => DATA <= x"FD";
            when x"5C7" => DATA <= x"FE";
            when x"5C8" => DATA <= x"2C";
            when x"5C9" => DATA <= x"FD";
            when x"5CA" => DATA <= x"FE";
            when x"5CB" => DATA <= x"2C";
            when x"5CC" => DATA <= x"FE";
            when x"5CD" => DATA <= x"FE";
            when x"5CE" => DATA <= x"10";
            when x"5CF" => DATA <= x"FB";
            when x"5D0" => DATA <= x"AD";
            when x"5D1" => DATA <= x"FF";
            when x"5D2" => DATA <= x"FE";
            when x"5D3" => DATA <= x"68";
            when x"5D4" => DATA <= x"C9";
            when x"5D5" => DATA <= x"06";
            when x"5D6" => DATA <= x"90";
            when x"5D7" => DATA <= x"1C";
            when x"5D8" => DATA <= x"D0";
            when x"5D9" => DATA <= x"1F";
            when x"5DA" => DATA <= x"A0";
            when x"5DB" => DATA <= x"00";
            when x"5DC" => DATA <= x"AD";
            when x"5DD" => DATA <= x"FC";
            when x"5DE" => DATA <= x"FE";
            when x"5DF" => DATA <= x"29";
            when x"5E0" => DATA <= x"80";
            when x"5E1" => DATA <= x"10";
            when x"5E2" => DATA <= x"F9";
            when x"5E3" => DATA <= x"B9";
            when x"5E4" => DATA <= x"FF";
            when x"5E5" => DATA <= x"FF";
            when x"5E6" => DATA <= x"8D";
            when x"5E7" => DATA <= x"FD";
            when x"5E8" => DATA <= x"FE";
            when x"5E9" => DATA <= x"C8";
            when x"5EA" => DATA <= x"D0";
            when x"5EB" => DATA <= x"F0";
            when x"5EC" => DATA <= x"2C";
            when x"5ED" => DATA <= x"FC";
            when x"5EE" => DATA <= x"FE";
            when x"5EF" => DATA <= x"10";
            when x"5F0" => DATA <= x"FB";
            when x"5F1" => DATA <= x"8D";
            when x"5F2" => DATA <= x"FD";
            when x"5F3" => DATA <= x"FE";
            when x"5F4" => DATA <= x"68";
            when x"5F5" => DATA <= x"A8";
            when x"5F6" => DATA <= x"A5";
            when x"5F7" => DATA <= x"FC";
            when x"5F8" => DATA <= x"40";
            when x"5F9" => DATA <= x"A0";
            when x"5FA" => DATA <= x"00";
            when x"5FB" => DATA <= x"AD";
            when x"5FC" => DATA <= x"FC";
            when x"5FD" => DATA <= x"FE";
            when x"5FE" => DATA <= x"29";
            when x"5FF" => DATA <= x"80";
            when x"600" => DATA <= x"10";
            when x"601" => DATA <= x"F9";
            when x"602" => DATA <= x"AD";
            when x"603" => DATA <= x"FD";
            when x"604" => DATA <= x"FE";
            when x"605" => DATA <= x"99";
            when x"606" => DATA <= x"FF";
            when x"607" => DATA <= x"FF";
            when x"608" => DATA <= x"C8";
            when x"609" => DATA <= x"D0";
            when x"60A" => DATA <= x"F0";
            when x"60B" => DATA <= x"F0";
            when x"60C" => DATA <= x"E7";
            when x"60D" => DATA <= x"48";
            when x"60E" => DATA <= x"AD";
            when x"60F" => DATA <= x"FF";
            when x"610" => DATA <= x"FF";
            when x"611" => DATA <= x"8D";
            when x"612" => DATA <= x"FD";
            when x"613" => DATA <= x"FE";
            when x"614" => DATA <= x"EE";
            when x"615" => DATA <= x"0F";
            when x"616" => DATA <= x"FE";
            when x"617" => DATA <= x"D0";
            when x"618" => DATA <= x"03";
            when x"619" => DATA <= x"EE";
            when x"61A" => DATA <= x"10";
            when x"61B" => DATA <= x"FE";
            when x"61C" => DATA <= x"68";
            when x"61D" => DATA <= x"40";
            when x"61E" => DATA <= x"48";
            when x"61F" => DATA <= x"AD";
            when x"620" => DATA <= x"FD";
            when x"621" => DATA <= x"FE";
            when x"622" => DATA <= x"8D";
            when x"623" => DATA <= x"FF";
            when x"624" => DATA <= x"FF";
            when x"625" => DATA <= x"EE";
            when x"626" => DATA <= x"23";
            when x"627" => DATA <= x"FE";
            when x"628" => DATA <= x"D0";
            when x"629" => DATA <= x"03";
            when x"62A" => DATA <= x"EE";
            when x"62B" => DATA <= x"24";
            when x"62C" => DATA <= x"FE";
            when x"62D" => DATA <= x"68";
            when x"62E" => DATA <= x"40";
            when x"62F" => DATA <= x"48";
            when x"630" => DATA <= x"98";
            when x"631" => DATA <= x"48";
            when x"632" => DATA <= x"A0";
            when x"633" => DATA <= x"00";
            when x"634" => DATA <= x"B1";
            when x"635" => DATA <= x"F6";
            when x"636" => DATA <= x"8D";
            when x"637" => DATA <= x"FD";
            when x"638" => DATA <= x"FE";
            when x"639" => DATA <= x"E6";
            when x"63A" => DATA <= x"F6";
            when x"63B" => DATA <= x"D0";
            when x"63C" => DATA <= x"02";
            when x"63D" => DATA <= x"E6";
            when x"63E" => DATA <= x"F7";
            when x"63F" => DATA <= x"B1";
            when x"640" => DATA <= x"F6";
            when x"641" => DATA <= x"8D";
            when x"642" => DATA <= x"FD";
            when x"643" => DATA <= x"FE";
            when x"644" => DATA <= x"E6";
            when x"645" => DATA <= x"F6";
            when x"646" => DATA <= x"D0";
            when x"647" => DATA <= x"02";
            when x"648" => DATA <= x"E6";
            when x"649" => DATA <= x"F7";
            when x"64A" => DATA <= x"68";
            when x"64B" => DATA <= x"A8";
            when x"64C" => DATA <= x"68";
            when x"64D" => DATA <= x"40";
            when x"64E" => DATA <= x"48";
            when x"64F" => DATA <= x"98";
            when x"650" => DATA <= x"48";
            when x"651" => DATA <= x"A0";
            when x"652" => DATA <= x"00";
            when x"653" => DATA <= x"AD";
            when x"654" => DATA <= x"FD";
            when x"655" => DATA <= x"FE";
            when x"656" => DATA <= x"91";
            when x"657" => DATA <= x"F6";
            when x"658" => DATA <= x"E6";
            when x"659" => DATA <= x"F6";
            when x"65A" => DATA <= x"D0";
            when x"65B" => DATA <= x"02";
            when x"65C" => DATA <= x"E6";
            when x"65D" => DATA <= x"F7";
            when x"65E" => DATA <= x"AD";
            when x"65F" => DATA <= x"FD";
            when x"660" => DATA <= x"FE";
            when x"661" => DATA <= x"91";
            when x"662" => DATA <= x"F6";
            when x"663" => DATA <= x"E6";
            when x"664" => DATA <= x"F6";
            when x"665" => DATA <= x"D0";
            when x"666" => DATA <= x"02";
            when x"667" => DATA <= x"E6";
            when x"668" => DATA <= x"F7";
            when x"669" => DATA <= x"68";
            when x"66A" => DATA <= x"A8";
            when x"66B" => DATA <= x"68";
            when x"66C" => DATA <= x"40";
            when x"66D" => DATA <= x"0F";
            when x"66E" => DATA <= x"23";
            when x"66F" => DATA <= x"F6";
            when x"670" => DATA <= x"F6";
            when x"671" => DATA <= x"F6";
            when x"672" => DATA <= x"F6";
            when x"673" => DATA <= x"E4";
            when x"674" => DATA <= x"06";
            when x"675" => DATA <= x"FE";
            when x"676" => DATA <= x"FE";
            when x"677" => DATA <= x"00";
            when x"678" => DATA <= x"00";
            when x"679" => DATA <= x"00";
            when x"67A" => DATA <= x"00";
            when x"67B" => DATA <= x"FD";
            when x"67C" => DATA <= x"FE";
            when x"67D" => DATA <= x"0D";
            when x"67E" => DATA <= x"1E";
            when x"67F" => DATA <= x"2F";
            when x"680" => DATA <= x"4E";
            when x"681" => DATA <= x"C0";
            when x"682" => DATA <= x"C0";
            when x"683" => DATA <= x"C0";
            when x"684" => DATA <= x"C0";
            when x"685" => DATA <= x"FE";
            when x"686" => DATA <= x"FE";
            when x"687" => DATA <= x"FE";
            when x"688" => DATA <= x"FE";
            when x"689" => DATA <= x"FE";
            when x"68A" => DATA <= x"FE";
            when x"68B" => DATA <= x"FE";
            when x"68C" => DATA <= x"FE";
            when x"68D" => DATA <= x"2C";
            when x"68E" => DATA <= x"F8";
            when x"68F" => DATA <= x"FE";
            when x"690" => DATA <= x"30";
            when x"691" => DATA <= x"0F";
            when x"692" => DATA <= x"2C";
            when x"693" => DATA <= x"FE";
            when x"694" => DATA <= x"FE";
            when x"695" => DATA <= x"10";
            when x"696" => DATA <= x"F6";
            when x"697" => DATA <= x"A5";
            when x"698" => DATA <= x"FC";
            when x"699" => DATA <= x"08";
            when x"69A" => DATA <= x"58";
            when x"69B" => DATA <= x"28";
            when x"69C" => DATA <= x"85";
            when x"69D" => DATA <= x"FC";
            when x"69E" => DATA <= x"4C";
            when x"69F" => DATA <= x"8D";
            when x"6A0" => DATA <= x"FE";
            when x"6A1" => DATA <= x"AD";
            when x"6A2" => DATA <= x"F9";
            when x"6A3" => DATA <= x"FE";
            when x"6A4" => DATA <= x"60";
            when x"6A5" => DATA <= x"68";
            when x"6A6" => DATA <= x"85";
            when x"6A7" => DATA <= x"FA";
            when x"6A8" => DATA <= x"68";
            when x"6A9" => DATA <= x"85";
            when x"6AA" => DATA <= x"FB";
            when x"6AB" => DATA <= x"A0";
            when x"6AC" => DATA <= x"00";
            when x"6AD" => DATA <= x"E6";
            when x"6AE" => DATA <= x"FA";
            when x"6AF" => DATA <= x"D0";
            when x"6B0" => DATA <= x"02";
            when x"6B1" => DATA <= x"E6";
            when x"6B2" => DATA <= x"FB";
            when x"6B3" => DATA <= x"B1";
            when x"6B4" => DATA <= x"FA";
            when x"6B5" => DATA <= x"30";
            when x"6B6" => DATA <= x"06";
            when x"6B7" => DATA <= x"20";
            when x"6B8" => DATA <= x"EE";
            when x"6B9" => DATA <= x"FF";
            when x"6BA" => DATA <= x"4C";
            when x"6BB" => DATA <= x"AD";
            when x"6BC" => DATA <= x"FE";
            when x"6BD" => DATA <= x"6C";
            when x"6BE" => DATA <= x"FA";
            when x"6BF" => DATA <= x"00";
            when x"6C0" => DATA <= x"8D";
            when x"6C1" => DATA <= x"FD";
            when x"6C2" => DATA <= x"FE";
            when x"6C3" => DATA <= x"40";
            when x"6C4" => DATA <= x"FF";
            when x"6C5" => DATA <= x"FF";
            when x"6C6" => DATA <= x"FF";
            when x"6C7" => DATA <= x"FF";
            when x"6C8" => DATA <= x"FF";
            when x"6C9" => DATA <= x"FF";
            when x"6CA" => DATA <= x"FF";
            when x"6CB" => DATA <= x"FF";
            when x"6CC" => DATA <= x"FF";
            when x"6CD" => DATA <= x"FF";
            when x"6CE" => DATA <= x"FF";
            when x"6CF" => DATA <= x"FF";
            when x"6D0" => DATA <= x"FF";
            when x"6D1" => DATA <= x"FF";
            when x"6D2" => DATA <= x"FF";
            when x"6D3" => DATA <= x"FF";
            when x"6D4" => DATA <= x"FF";
            when x"6D5" => DATA <= x"FF";
            when x"6D6" => DATA <= x"FF";
            when x"6D7" => DATA <= x"FF";
            when x"6D8" => DATA <= x"FF";
            when x"6D9" => DATA <= x"FF";
            when x"6DA" => DATA <= x"FF";
            when x"6DB" => DATA <= x"FF";
            when x"6DC" => DATA <= x"FF";
            when x"6DD" => DATA <= x"FF";
            when x"6DE" => DATA <= x"FF";
            when x"6DF" => DATA <= x"FF";
            when x"6E0" => DATA <= x"FF";
            when x"6E1" => DATA <= x"FF";
            when x"6E2" => DATA <= x"FF";
            when x"6E3" => DATA <= x"FF";
            when x"6E4" => DATA <= x"FF";
            when x"6E5" => DATA <= x"FF";
            when x"6E6" => DATA <= x"FF";
            when x"6E7" => DATA <= x"FF";
            when x"6E8" => DATA <= x"FF";
            when x"6E9" => DATA <= x"FF";
            when x"6EA" => DATA <= x"FF";
            when x"6EB" => DATA <= x"FF";
            when x"6EC" => DATA <= x"FF";
            when x"6ED" => DATA <= x"FF";
            when x"6EE" => DATA <= x"FF";
            when x"6EF" => DATA <= x"FF";
            when x"6F0" => DATA <= x"00";
            when x"6F1" => DATA <= x"00";
            when x"6F2" => DATA <= x"00";
            when x"6F3" => DATA <= x"00";
            when x"6F4" => DATA <= x"00";
            when x"6F5" => DATA <= x"00";
            when x"6F6" => DATA <= x"00";
            when x"6F7" => DATA <= x"00";
            when x"6F8" => DATA <= x"00";
            when x"6F9" => DATA <= x"00";
            when x"6FA" => DATA <= x"00";
            when x"6FB" => DATA <= x"00";
            when x"6FC" => DATA <= x"00";
            when x"6FD" => DATA <= x"00";
            when x"6FE" => DATA <= x"00";
            when x"6FF" => DATA <= x"00";
            when x"700" => DATA <= x"FF";
            when x"701" => DATA <= x"FF";
            when x"702" => DATA <= x"FF";
            when x"703" => DATA <= x"FF";
            when x"704" => DATA <= x"FF";
            when x"705" => DATA <= x"FF";
            when x"706" => DATA <= x"FF";
            when x"707" => DATA <= x"FF";
            when x"708" => DATA <= x"FF";
            when x"709" => DATA <= x"FF";
            when x"70A" => DATA <= x"FF";
            when x"70B" => DATA <= x"FF";
            when x"70C" => DATA <= x"FF";
            when x"70D" => DATA <= x"FF";
            when x"70E" => DATA <= x"FF";
            when x"70F" => DATA <= x"FF";
            when x"710" => DATA <= x"FF";
            when x"711" => DATA <= x"FF";
            when x"712" => DATA <= x"FF";
            when x"713" => DATA <= x"FF";
            when x"714" => DATA <= x"FF";
            when x"715" => DATA <= x"FF";
            when x"716" => DATA <= x"FF";
            when x"717" => DATA <= x"FF";
            when x"718" => DATA <= x"FF";
            when x"719" => DATA <= x"FF";
            when x"71A" => DATA <= x"FF";
            when x"71B" => DATA <= x"FF";
            when x"71C" => DATA <= x"FF";
            when x"71D" => DATA <= x"FF";
            when x"71E" => DATA <= x"FF";
            when x"71F" => DATA <= x"FF";
            when x"720" => DATA <= x"FF";
            when x"721" => DATA <= x"FF";
            when x"722" => DATA <= x"FF";
            when x"723" => DATA <= x"FF";
            when x"724" => DATA <= x"FF";
            when x"725" => DATA <= x"FF";
            when x"726" => DATA <= x"FF";
            when x"727" => DATA <= x"FF";
            when x"728" => DATA <= x"FF";
            when x"729" => DATA <= x"FF";
            when x"72A" => DATA <= x"FF";
            when x"72B" => DATA <= x"FF";
            when x"72C" => DATA <= x"FF";
            when x"72D" => DATA <= x"FF";
            when x"72E" => DATA <= x"FF";
            when x"72F" => DATA <= x"FF";
            when x"730" => DATA <= x"FF";
            when x"731" => DATA <= x"FF";
            when x"732" => DATA <= x"FF";
            when x"733" => DATA <= x"FF";
            when x"734" => DATA <= x"FF";
            when x"735" => DATA <= x"FF";
            when x"736" => DATA <= x"FF";
            when x"737" => DATA <= x"FF";
            when x"738" => DATA <= x"FF";
            when x"739" => DATA <= x"FF";
            when x"73A" => DATA <= x"FF";
            when x"73B" => DATA <= x"FF";
            when x"73C" => DATA <= x"FF";
            when x"73D" => DATA <= x"FF";
            when x"73E" => DATA <= x"FF";
            when x"73F" => DATA <= x"FF";
            when x"740" => DATA <= x"FF";
            when x"741" => DATA <= x"FF";
            when x"742" => DATA <= x"FF";
            when x"743" => DATA <= x"FF";
            when x"744" => DATA <= x"FF";
            when x"745" => DATA <= x"FF";
            when x"746" => DATA <= x"FF";
            when x"747" => DATA <= x"FF";
            when x"748" => DATA <= x"FF";
            when x"749" => DATA <= x"FF";
            when x"74A" => DATA <= x"FF";
            when x"74B" => DATA <= x"FF";
            when x"74C" => DATA <= x"FF";
            when x"74D" => DATA <= x"FF";
            when x"74E" => DATA <= x"FF";
            when x"74F" => DATA <= x"FF";
            when x"750" => DATA <= x"FF";
            when x"751" => DATA <= x"FF";
            when x"752" => DATA <= x"FF";
            when x"753" => DATA <= x"FF";
            when x"754" => DATA <= x"FF";
            when x"755" => DATA <= x"FF";
            when x"756" => DATA <= x"FF";
            when x"757" => DATA <= x"FF";
            when x"758" => DATA <= x"FF";
            when x"759" => DATA <= x"FF";
            when x"75A" => DATA <= x"FF";
            when x"75B" => DATA <= x"FF";
            when x"75C" => DATA <= x"FF";
            when x"75D" => DATA <= x"FF";
            when x"75E" => DATA <= x"FF";
            when x"75F" => DATA <= x"FF";
            when x"760" => DATA <= x"FF";
            when x"761" => DATA <= x"FF";
            when x"762" => DATA <= x"FF";
            when x"763" => DATA <= x"FF";
            when x"764" => DATA <= x"FF";
            when x"765" => DATA <= x"FF";
            when x"766" => DATA <= x"FF";
            when x"767" => DATA <= x"FF";
            when x"768" => DATA <= x"FF";
            when x"769" => DATA <= x"FF";
            when x"76A" => DATA <= x"FF";
            when x"76B" => DATA <= x"FF";
            when x"76C" => DATA <= x"FF";
            when x"76D" => DATA <= x"FF";
            when x"76E" => DATA <= x"FF";
            when x"76F" => DATA <= x"FF";
            when x"770" => DATA <= x"FF";
            when x"771" => DATA <= x"FF";
            when x"772" => DATA <= x"FF";
            when x"773" => DATA <= x"FF";
            when x"774" => DATA <= x"FF";
            when x"775" => DATA <= x"FF";
            when x"776" => DATA <= x"FF";
            when x"777" => DATA <= x"FF";
            when x"778" => DATA <= x"FF";
            when x"779" => DATA <= x"FF";
            when x"77A" => DATA <= x"FF";
            when x"77B" => DATA <= x"FF";
            when x"77C" => DATA <= x"FF";
            when x"77D" => DATA <= x"FF";
            when x"77E" => DATA <= x"FF";
            when x"77F" => DATA <= x"FF";
            when x"780" => DATA <= x"C4";
            when x"781" => DATA <= x"FC";
            when x"782" => DATA <= x"50";
            when x"783" => DATA <= x"F9";
            when x"784" => DATA <= x"FD";
            when x"785" => DATA <= x"FC";
            when x"786" => DATA <= x"C4";
            when x"787" => DATA <= x"FC";
            when x"788" => DATA <= x"D5";
            when x"789" => DATA <= x"F9";
            when x"78A" => DATA <= x"80";
            when x"78B" => DATA <= x"FA";
            when x"78C" => DATA <= x"0C";
            when x"78D" => DATA <= x"FB";
            when x"78E" => DATA <= x"6D";
            when x"78F" => DATA <= x"F9";
            when x"790" => DATA <= x"77";
            when x"791" => DATA <= x"F9";
            when x"792" => DATA <= x"60";
            when x"793" => DATA <= x"FC";
            when x"794" => DATA <= x"D9";
            when x"795" => DATA <= x"FB";
            when x"796" => DATA <= x"37";
            when x"797" => DATA <= x"FC";
            when x"798" => DATA <= x"43";
            when x"799" => DATA <= x"FC";
            when x"79A" => DATA <= x"9B";
            when x"79B" => DATA <= x"FC";
            when x"79C" => DATA <= x"19";
            when x"79D" => DATA <= x"FC";
            when x"79E" => DATA <= x"C4";
            when x"79F" => DATA <= x"FC";
            when x"7A0" => DATA <= x"88";
            when x"7A1" => DATA <= x"F9";
            when x"7A2" => DATA <= x"C4";
            when x"7A3" => DATA <= x"FC";
            when x"7A4" => DATA <= x"C4";
            when x"7A5" => DATA <= x"FC";
            when x"7A6" => DATA <= x"C4";
            when x"7A7" => DATA <= x"FC";
            when x"7A8" => DATA <= x"C4";
            when x"7A9" => DATA <= x"FC";
            when x"7AA" => DATA <= x"C4";
            when x"7AB" => DATA <= x"FC";
            when x"7AC" => DATA <= x"C4";
            when x"7AD" => DATA <= x"FC";
            when x"7AE" => DATA <= x"C4";
            when x"7AF" => DATA <= x"FC";
            when x"7B0" => DATA <= x"88";
            when x"7B1" => DATA <= x"F9";
            when x"7B2" => DATA <= x"88";
            when x"7B3" => DATA <= x"F9";
            when x"7B4" => DATA <= x"88";
            when x"7B5" => DATA <= x"F9";
            when x"7B6" => DATA <= x"36";
            when x"7B7" => DATA <= x"80";
            when x"7B8" => DATA <= x"FF";
            when x"7B9" => DATA <= x"4C";
            when x"7BA" => DATA <= x"C4";
            when x"7BB" => DATA <= x"FC";
            when x"7BC" => DATA <= x"4C";
            when x"7BD" => DATA <= x"C4";
            when x"7BE" => DATA <= x"FC";
            when x"7BF" => DATA <= x"4C";
            when x"7C0" => DATA <= x"C4";
            when x"7C1" => DATA <= x"FC";
            when x"7C2" => DATA <= x"4C";
            when x"7C3" => DATA <= x"C4";
            when x"7C4" => DATA <= x"FC";
            when x"7C5" => DATA <= x"4C";
            when x"7C6" => DATA <= x"C4";
            when x"7C7" => DATA <= x"FC";
            when x"7C8" => DATA <= x"4C";
            when x"7C9" => DATA <= x"77";
            when x"7CA" => DATA <= x"F9";
            when x"7CB" => DATA <= x"4C";
            when x"7CC" => DATA <= x"6D";
            when x"7CD" => DATA <= x"F9";
            when x"7CE" => DATA <= x"6C";
            when x"7CF" => DATA <= x"1C";
            when x"7D0" => DATA <= x"02";
            when x"7D1" => DATA <= x"6C";
            when x"7D2" => DATA <= x"1A";
            when x"7D3" => DATA <= x"02";
            when x"7D4" => DATA <= x"6C";
            when x"7D5" => DATA <= x"18";
            when x"7D6" => DATA <= x"02";
            when x"7D7" => DATA <= x"6C";
            when x"7D8" => DATA <= x"16";
            when x"7D9" => DATA <= x"02";
            when x"7DA" => DATA <= x"6C";
            when x"7DB" => DATA <= x"14";
            when x"7DC" => DATA <= x"02";
            when x"7DD" => DATA <= x"6C";
            when x"7DE" => DATA <= x"12";
            when x"7DF" => DATA <= x"02";
            when x"7E0" => DATA <= x"6C";
            when x"7E1" => DATA <= x"10";
            when x"7E2" => DATA <= x"02";
            when x"7E3" => DATA <= x"C9";
            when x"7E4" => DATA <= x"0D";
            when x"7E5" => DATA <= x"D0";
            when x"7E6" => DATA <= x"07";
            when x"7E7" => DATA <= x"A9";
            when x"7E8" => DATA <= x"0A";
            when x"7E9" => DATA <= x"20";
            when x"7EA" => DATA <= x"EE";
            when x"7EB" => DATA <= x"FF";
            when x"7EC" => DATA <= x"A9";
            when x"7ED" => DATA <= x"0D";
            when x"7EE" => DATA <= x"6C";
            when x"7EF" => DATA <= x"0E";
            when x"7F0" => DATA <= x"02";
            when x"7F1" => DATA <= x"6C";
            when x"7F2" => DATA <= x"0C";
            when x"7F3" => DATA <= x"02";
            when x"7F4" => DATA <= x"6C";
            when x"7F5" => DATA <= x"0A";
            when x"7F6" => DATA <= x"02";
            when x"7F7" => DATA <= x"6C";
            when x"7F8" => DATA <= x"08";
            when x"7F9" => DATA <= x"02";
            when x"7FA" => DATA <= x"0D";
            when x"7FB" => DATA <= x"FE";
            when x"7FC" => DATA <= x"00";
            when x"7FD" => DATA <= x"F8";
            when x"7FE" => DATA <= x"F2";
            when x"7FF" => DATA <= x"FC";
            when others => DATA <= (others => '0');
        end case;
    end process;
end RTL;
