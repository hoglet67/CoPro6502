library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tuberom_6809 is
    port (
        CLK  : in  std_logic;
        ADDR : in  std_logic_vector(10 downto 0);
        DATA : out std_logic_vector(7 downto 0)
        );
end;

architecture RTL of tuberom_6809 is

    signal rom_addr : std_logic_vector(11 downto 0);

begin

    p_addr : process(ADDR)
    begin
        rom_addr              <= (others => '0');
        rom_addr(10 downto 0) <= ADDR;
    end process;

    p_rom : process
    begin
        wait until rising_edge(CLK);
        DATA <= (others => '0');
        case rom_addr is
            when x"000" => DATA <= x"F8";
            when x"001" => DATA <= x"2D";
            when x"002" => DATA <= x"F8";
            when x"003" => DATA <= x"67";
            when x"004" => DATA <= x"FF";
            when x"005" => DATA <= x"E0";
            when x"006" => DATA <= x"F8";
            when x"007" => DATA <= x"D0";
            when x"008" => DATA <= x"F8";
            when x"009" => DATA <= x"E4";
            when x"00A" => DATA <= x"FF";
            when x"00B" => DATA <= x"EE";
            when x"00C" => DATA <= x"F8";
            when x"00D" => DATA <= x"D9";
            when x"00E" => DATA <= x"FF";
            when x"00F" => DATA <= x"E7";
            when x"010" => DATA <= x"F8";
            when x"011" => DATA <= x"D6";
            when x"012" => DATA <= x"F8";
            when x"013" => DATA <= x"CF";
            when x"014" => DATA <= x"20";
            when x"015" => DATA <= x"51";
            when x"016" => DATA <= x"0D";
            when x"017" => DATA <= x"36";
            when x"018" => DATA <= x"38";
            when x"019" => DATA <= x"30";
            when x"01A" => DATA <= x"39";
            when x"01B" => DATA <= x"20";
            when x"01C" => DATA <= x"54";
            when x"01D" => DATA <= x"55";
            when x"01E" => DATA <= x"42";
            when x"01F" => DATA <= x"45";
            when x"020" => DATA <= x"20";
            when x"021" => DATA <= x"36";
            when x"022" => DATA <= x"34";
            when x"023" => DATA <= x"4B";
            when x"024" => DATA <= x"20";
            when x"025" => DATA <= x"76";
            when x"026" => DATA <= x"30";
            when x"027" => DATA <= x"2E";
            when x"028" => DATA <= x"32";
            when x"029" => DATA <= x"33";
            when x"02A" => DATA <= x"0D";
            when x"02B" => DATA <= x"0D";
            when x"02C" => DATA <= x"00";
            when x"02D" => DATA <= x"1A";
            when x"02E" => DATA <= x"50";
            when x"02F" => DATA <= x"10";
            when x"030" => DATA <= x"CE";
            when x"031" => DATA <= x"F8";
            when x"032" => DATA <= x"00";
            when x"033" => DATA <= x"1F";
            when x"034" => DATA <= x"41";
            when x"035" => DATA <= x"A6";
            when x"036" => DATA <= x"84";
            when x"037" => DATA <= x"A7";
            when x"038" => DATA <= x"80";
            when x"039" => DATA <= x"8C";
            when x"03A" => DATA <= x"FE";
            when x"03B" => DATA <= x"C0";
            when x"03C" => DATA <= x"26";
            when x"03D" => DATA <= x"F7";
            when x"03E" => DATA <= x"8E";
            when x"03F" => DATA <= x"FE";
            when x"040" => DATA <= x"F0";
            when x"041" => DATA <= x"A6";
            when x"042" => DATA <= x"84";
            when x"043" => DATA <= x"A7";
            when x"044" => DATA <= x"80";
            when x"045" => DATA <= x"8C";
            when x"046" => DATA <= x"00";
            when x"047" => DATA <= x"00";
            when x"048" => DATA <= x"26";
            when x"049" => DATA <= x"F7";
            when x"04A" => DATA <= x"B6";
            when x"04B" => DATA <= x"FE";
            when x"04C" => DATA <= x"E0";
            when x"04D" => DATA <= x"1A";
            when x"04E" => DATA <= x"50";
            when x"04F" => DATA <= x"10";
            when x"050" => DATA <= x"CE";
            when x"051" => DATA <= x"FF";
            when x"052" => DATA <= x"20";
            when x"053" => DATA <= x"BD";
            when x"054" => DATA <= x"F8";
            when x"055" => DATA <= x"B7";
            when x"056" => DATA <= x"1C";
            when x"057" => DATA <= x"00";
            when x"058" => DATA <= x"8E";
            when x"059" => DATA <= x"F8";
            when x"05A" => DATA <= x"16";
            when x"05B" => DATA <= x"BD";
            when x"05C" => DATA <= x"F9";
            when x"05D" => DATA <= x"24";
            when x"05E" => DATA <= x"B7";
            when x"05F" => DATA <= x"FF";
            when x"060" => DATA <= x"80";
            when x"061" => DATA <= x"BD";
            when x"062" => DATA <= x"FF";
            when x"063" => DATA <= x"EE";
            when x"064" => DATA <= x"BD";
            when x"065" => DATA <= x"F9";
            when x"066" => DATA <= x"56";
            when x"067" => DATA <= x"10";
            when x"068" => DATA <= x"CE";
            when x"069" => DATA <= x"FF";
            when x"06A" => DATA <= x"20";
            when x"06B" => DATA <= x"BD";
            when x"06C" => DATA <= x"F8";
            when x"06D" => DATA <= x"B7";
            when x"06E" => DATA <= x"10";
            when x"06F" => DATA <= x"FE";
            when x"070" => DATA <= x"FF";
            when x"071" => DATA <= x"8A";
            when x"072" => DATA <= x"1C";
            when x"073" => DATA <= x"00";
            when x"074" => DATA <= x"8E";
            when x"075" => DATA <= x"F8";
            when x"076" => DATA <= x"87";
            when x"077" => DATA <= x"BD";
            when x"078" => DATA <= x"F9";
            when x"079" => DATA <= x"24";
            when x"07A" => DATA <= x"BD";
            when x"07B" => DATA <= x"FF";
            when x"07C" => DATA <= x"F1";
            when x"07D" => DATA <= x"25";
            when x"07E" => DATA <= x"1D";
            when x"07F" => DATA <= x"8E";
            when x"080" => DATA <= x"FF";
            when x"081" => DATA <= x"20";
            when x"082" => DATA <= x"BD";
            when x"083" => DATA <= x"FF";
            when x"084" => DATA <= x"F7";
            when x"085" => DATA <= x"20";
            when x"086" => DATA <= x"E0";
            when x"087" => DATA <= x"36";
            when x"088" => DATA <= x"38";
            when x"089" => DATA <= x"30";
            when x"08A" => DATA <= x"39";
            when x"08B" => DATA <= x"3E";
            when x"08C" => DATA <= x"2A";
            when x"08D" => DATA <= x"00";
            when x"08E" => DATA <= x"FF";
            when x"08F" => DATA <= x"20";
            when x"090" => DATA <= x"5F";
            when x"091" => DATA <= x"20";
            when x"092" => DATA <= x"FF";
            when x"093" => DATA <= x"3F";
            when x"094" => DATA <= x"11";
            when x"095" => DATA <= x"45";
            when x"096" => DATA <= x"73";
            when x"097" => DATA <= x"63";
            when x"098" => DATA <= x"61";
            when x"099" => DATA <= x"70";
            when x"09A" => DATA <= x"65";
            when x"09B" => DATA <= x"00";
            when x"09C" => DATA <= x"86";
            when x"09D" => DATA <= x"7C";
            when x"09E" => DATA <= x"BD";
            when x"09F" => DATA <= x"FF";
            when x"0A0" => DATA <= x"F4";
            when x"0A1" => DATA <= x"8E";
            when x"0A2" => DATA <= x"F8";
            when x"0A3" => DATA <= x"94";
            when x"0A4" => DATA <= x"7E";
            when x"0A5" => DATA <= x"FF";
            when x"0A6" => DATA <= x"BC";
            when x"0A7" => DATA <= x"10";
            when x"0A8" => DATA <= x"FE";
            when x"0A9" => DATA <= x"FF";
            when x"0AA" => DATA <= x"8A";
            when x"0AB" => DATA <= x"BD";
            when x"0AC" => DATA <= x"FF";
            when x"0AD" => DATA <= x"E7";
            when x"0AE" => DATA <= x"A6";
            when x"0AF" => DATA <= x"80";
            when x"0B0" => DATA <= x"8D";
            when x"0B1" => DATA <= x"72";
            when x"0B2" => DATA <= x"BD";
            when x"0B3" => DATA <= x"FF";
            when x"0B4" => DATA <= x"E7";
            when x"0B5" => DATA <= x"20";
            when x"0B6" => DATA <= x"B0";
            when x"0B7" => DATA <= x"CC";
            when x"0B8" => DATA <= x"00";
            when x"0B9" => DATA <= x"00";
            when x"0BA" => DATA <= x"FD";
            when x"0BB" => DATA <= x"FF";
            when x"0BC" => DATA <= x"88";
            when x"0BD" => DATA <= x"CC";
            when x"0BE" => DATA <= x"F8";
            when x"0BF" => DATA <= x"00";
            when x"0C0" => DATA <= x"FD";
            when x"0C1" => DATA <= x"FF";
            when x"0C2" => DATA <= x"8A";
            when x"0C3" => DATA <= x"CC";
            when x"0C4" => DATA <= x"FD";
            when x"0C5" => DATA <= x"3D";
            when x"0C6" => DATA <= x"FD";
            when x"0C7" => DATA <= x"FE";
            when x"0C8" => DATA <= x"FA";
            when x"0C9" => DATA <= x"CC";
            when x"0CA" => DATA <= x"F8";
            when x"0CB" => DATA <= x"A7";
            when x"0CC" => DATA <= x"FD";
            when x"0CD" => DATA <= x"FF";
            when x"0CE" => DATA <= x"FA";
            when x"0CF" => DATA <= x"39";
            when x"0D0" => DATA <= x"BD";
            when x"0D1" => DATA <= x"FF";
            when x"0D2" => DATA <= x"E0";
            when x"0D3" => DATA <= x"7E";
            when x"0D4" => DATA <= x"FF";
            when x"0D5" => DATA <= x"EE";
            when x"0D6" => DATA <= x"BD";
            when x"0D7" => DATA <= x"FF";
            when x"0D8" => DATA <= x"E7";
            when x"0D9" => DATA <= x"A6";
            when x"0DA" => DATA <= x"80";
            when x"0DB" => DATA <= x"81";
            when x"0DC" => DATA <= x"04";
            when x"0DD" => DATA <= x"27";
            when x"0DE" => DATA <= x"F0";
            when x"0DF" => DATA <= x"BD";
            when x"0E0" => DATA <= x"FF";
            when x"0E1" => DATA <= x"EE";
            when x"0E2" => DATA <= x"20";
            when x"0E3" => DATA <= x"F5";
            when x"0E4" => DATA <= x"34";
            when x"0E5" => DATA <= x"32";
            when x"0E6" => DATA <= x"86";
            when x"0E7" => DATA <= x"80";
            when x"0E8" => DATA <= x"8E";
            when x"0E9" => DATA <= x"FF";
            when x"0EA" => DATA <= x"FF";
            when x"0EB" => DATA <= x"1F";
            when x"0EC" => DATA <= x"12";
            when x"0ED" => DATA <= x"BD";
            when x"0EE" => DATA <= x"FF";
            when x"0EF" => DATA <= x"F4";
            when x"0F0" => DATA <= x"8C";
            when x"0F1" => DATA <= x"00";
            when x"0F2" => DATA <= x"00";
            when x"0F3" => DATA <= x"35";
            when x"0F4" => DATA <= x"B2";
            when x"0F5" => DATA <= x"34";
            when x"0F6" => DATA <= x"06";
            when x"0F7" => DATA <= x"1F";
            when x"0F8" => DATA <= x"10";
            when x"0F9" => DATA <= x"8D";
            when x"0FA" => DATA <= x"06";
            when x"0FB" => DATA <= x"1F";
            when x"0FC" => DATA <= x"98";
            when x"0FD" => DATA <= x"8D";
            when x"0FE" => DATA <= x"02";
            when x"0FF" => DATA <= x"35";
            when x"100" => DATA <= x"86";
            when x"101" => DATA <= x"34";
            when x"102" => DATA <= x"02";
            when x"103" => DATA <= x"44";
            when x"104" => DATA <= x"44";
            when x"105" => DATA <= x"44";
            when x"106" => DATA <= x"44";
            when x"107" => DATA <= x"8D";
            when x"108" => DATA <= x"06";
            when x"109" => DATA <= x"A6";
            when x"10A" => DATA <= x"E4";
            when x"10B" => DATA <= x"8D";
            when x"10C" => DATA <= x"02";
            when x"10D" => DATA <= x"35";
            when x"10E" => DATA <= x"82";
            when x"10F" => DATA <= x"84";
            when x"110" => DATA <= x"0F";
            when x"111" => DATA <= x"81";
            when x"112" => DATA <= x"0A";
            when x"113" => DATA <= x"25";
            when x"114" => DATA <= x"02";
            when x"115" => DATA <= x"8B";
            when x"116" => DATA <= x"07";
            when x"117" => DATA <= x"8B";
            when x"118" => DATA <= x"30";
            when x"119" => DATA <= x"7E";
            when x"11A" => DATA <= x"FF";
            when x"11B" => DATA <= x"EE";
            when x"11C" => DATA <= x"35";
            when x"11D" => DATA <= x"10";
            when x"11E" => DATA <= x"BD";
            when x"11F" => DATA <= x"F9";
            when x"120" => DATA <= x"24";
            when x"121" => DATA <= x"34";
            when x"122" => DATA <= x"10";
            when x"123" => DATA <= x"39";
            when x"124" => DATA <= x"A6";
            when x"125" => DATA <= x"80";
            when x"126" => DATA <= x"27";
            when x"127" => DATA <= x"FB";
            when x"128" => DATA <= x"BD";
            when x"129" => DATA <= x"FF";
            when x"12A" => DATA <= x"E3";
            when x"12B" => DATA <= x"20";
            when x"12C" => DATA <= x"F7";
            when x"12D" => DATA <= x"4F";
            when x"12E" => DATA <= x"BD";
            when x"12F" => DATA <= x"FB";
            when x"130" => DATA <= x"CA";
            when x"131" => DATA <= x"8D";
            when x"132" => DATA <= x"02";
            when x"133" => DATA <= x"8B";
            when x"134" => DATA <= x"80";
            when x"135" => DATA <= x"B6";
            when x"136" => DATA <= x"FE";
            when x"137" => DATA <= x"E2";
            when x"138" => DATA <= x"2A";
            when x"139" => DATA <= x"FB";
            when x"13A" => DATA <= x"B6";
            when x"13B" => DATA <= x"FE";
            when x"13C" => DATA <= x"E3";
            when x"13D" => DATA <= x"39";
            when x"13E" => DATA <= x"10";
            when x"13F" => DATA <= x"FF";
            when x"140" => DATA <= x"F9";
            when x"141" => DATA <= x"4B";
            when x"142" => DATA <= x"10";
            when x"143" => DATA <= x"CE";
            when x"144" => DATA <= x"FF";
            when x"145" => DATA <= x"20";
            when x"146" => DATA <= x"BD";
            when x"147" => DATA <= x"F9";
            when x"148" => DATA <= x"4E";
            when x"149" => DATA <= x"10";
            when x"14A" => DATA <= x"CE";
            when x"14B" => DATA <= x"00";
            when x"14C" => DATA <= x"00";
            when x"14D" => DATA <= x"39";
            when x"14E" => DATA <= x"86";
            when x"14F" => DATA <= x"02";
            when x"150" => DATA <= x"BD";
            when x"151" => DATA <= x"FB";
            when x"152" => DATA <= x"CA";
            when x"153" => DATA <= x"BD";
            when x"154" => DATA <= x"FB";
            when x"155" => DATA <= x"8F";
            when x"156" => DATA <= x"8D";
            when x"157" => DATA <= x"DD";
            when x"158" => DATA <= x"2A";
            when x"159" => DATA <= x"30";
            when x"15A" => DATA <= x"BE";
            when x"15B" => DATA <= x"FF";
            when x"15C" => DATA <= x"90";
            when x"15D" => DATA <= x"A6";
            when x"15E" => DATA <= x"07";
            when x"15F" => DATA <= x"A6";
            when x"160" => DATA <= x"86";
            when x"161" => DATA <= x"26";
            when x"162" => DATA <= x"0B";
            when x"163" => DATA <= x"A6";
            when x"164" => DATA <= x"06";
            when x"165" => DATA <= x"48";
            when x"166" => DATA <= x"2A";
            when x"167" => DATA <= x"23";
            when x"168" => DATA <= x"84";
            when x"169" => DATA <= x"1E";
            when x"16A" => DATA <= x"81";
            when x"16B" => DATA <= x"06";
            when x"16C" => DATA <= x"26";
            when x"16D" => DATA <= x"1D";
            when x"16E" => DATA <= x"10";
            when x"16F" => DATA <= x"BE";
            when x"170" => DATA <= x"FF";
            when x"171" => DATA <= x"8A";
            when x"172" => DATA <= x"34";
            when x"173" => DATA <= x"20";
            when x"174" => DATA <= x"8C";
            when x"175" => DATA <= x"80";
            when x"176" => DATA <= x"00";
            when x"177" => DATA <= x"25";
            when x"178" => DATA <= x"08";
            when x"179" => DATA <= x"8C";
            when x"17A" => DATA <= x"F8";
            when x"17B" => DATA <= x"00";
            when x"17C" => DATA <= x"24";
            when x"17D" => DATA <= x"03";
            when x"17E" => DATA <= x"BF";
            when x"17F" => DATA <= x"FF";
            when x"180" => DATA <= x"8A";
            when x"181" => DATA <= x"86";
            when x"182" => DATA <= x"01";
            when x"183" => DATA <= x"AD";
            when x"184" => DATA <= x"84";
            when x"185" => DATA <= x"35";
            when x"186" => DATA <= x"10";
            when x"187" => DATA <= x"BF";
            when x"188" => DATA <= x"FF";
            when x"189" => DATA <= x"8A";
            when x"18A" => DATA <= x"39";
            when x"18B" => DATA <= x"BD";
            when x"18C" => DATA <= x"FF";
            when x"18D" => DATA <= x"BF";
            when x"18E" => DATA <= x"3F";
            when x"18F" => DATA <= x"F7";
            when x"190" => DATA <= x"4E";
            when x"191" => DATA <= x"6F";
            when x"192" => DATA <= x"74";
            when x"193" => DATA <= x"20";
            when x"194" => DATA <= x"36";
            when x"195" => DATA <= x"38";
            when x"196" => DATA <= x"30";
            when x"197" => DATA <= x"39";
            when x"198" => DATA <= x"20";
            when x"199" => DATA <= x"63";
            when x"19A" => DATA <= x"6F";
            when x"19B" => DATA <= x"64";
            when x"19C" => DATA <= x"65";
            when x"19D" => DATA <= x"00";
            when x"19E" => DATA <= x"81";
            when x"19F" => DATA <= x"80";
            when x"1A0" => DATA <= x"24";
            when x"1A1" => DATA <= x"1D";
            when x"1A2" => DATA <= x"34";
            when x"1A3" => DATA <= x"06";
            when x"1A4" => DATA <= x"86";
            when x"1A5" => DATA <= x"04";
            when x"1A6" => DATA <= x"BD";
            when x"1A7" => DATA <= x"FB";
            when x"1A8" => DATA <= x"CA";
            when x"1A9" => DATA <= x"1F";
            when x"1AA" => DATA <= x"10";
            when x"1AB" => DATA <= x"BD";
            when x"1AC" => DATA <= x"FB";
            when x"1AD" => DATA <= x"C8";
            when x"1AE" => DATA <= x"35";
            when x"1AF" => DATA <= x"06";
            when x"1B0" => DATA <= x"34";
            when x"1B1" => DATA <= x"06";
            when x"1B2" => DATA <= x"BD";
            when x"1B3" => DATA <= x"FB";
            when x"1B4" => DATA <= x"CA";
            when x"1B5" => DATA <= x"BD";
            when x"1B6" => DATA <= x"F9";
            when x"1B7" => DATA <= x"35";
            when x"1B8" => DATA <= x"1F";
            when x"1B9" => DATA <= x"89";
            when x"1BA" => DATA <= x"4F";
            when x"1BB" => DATA <= x"1F";
            when x"1BC" => DATA <= x"01";
            when x"1BD" => DATA <= x"35";
            when x"1BE" => DATA <= x"86";
            when x"1BF" => DATA <= x"81";
            when x"1C0" => DATA <= x"82";
            when x"1C1" => DATA <= x"27";
            when x"1C2" => DATA <= x"42";
            when x"1C3" => DATA <= x"81";
            when x"1C4" => DATA <= x"83";
            when x"1C5" => DATA <= x"27";
            when x"1C6" => DATA <= x"42";
            when x"1C7" => DATA <= x"81";
            when x"1C8" => DATA <= x"84";
            when x"1C9" => DATA <= x"27";
            when x"1CA" => DATA <= x"42";
            when x"1CB" => DATA <= x"34";
            when x"1CC" => DATA <= x"06";
            when x"1CD" => DATA <= x"86";
            when x"1CE" => DATA <= x"06";
            when x"1CF" => DATA <= x"BD";
            when x"1D0" => DATA <= x"FB";
            when x"1D1" => DATA <= x"CA";
            when x"1D2" => DATA <= x"1F";
            when x"1D3" => DATA <= x"10";
            when x"1D4" => DATA <= x"BD";
            when x"1D5" => DATA <= x"FB";
            when x"1D6" => DATA <= x"C8";
            when x"1D7" => DATA <= x"1F";
            when x"1D8" => DATA <= x"20";
            when x"1D9" => DATA <= x"BD";
            when x"1DA" => DATA <= x"FB";
            when x"1DB" => DATA <= x"C8";
            when x"1DC" => DATA <= x"35";
            when x"1DD" => DATA <= x"06";
            when x"1DE" => DATA <= x"BD";
            when x"1DF" => DATA <= x"FB";
            when x"1E0" => DATA <= x"CA";
            when x"1E1" => DATA <= x"81";
            when x"1E2" => DATA <= x"9D";
            when x"1E3" => DATA <= x"27";
            when x"1E4" => DATA <= x"23";
            when x"1E5" => DATA <= x"81";
            when x"1E6" => DATA <= x"8E";
            when x"1E7" => DATA <= x"10";
            when x"1E8" => DATA <= x"27";
            when x"1E9" => DATA <= x"FF";
            when x"1EA" => DATA <= x"6B";
            when x"1EB" => DATA <= x"34";
            when x"1EC" => DATA <= x"06";
            when x"1ED" => DATA <= x"BD";
            when x"1EE" => DATA <= x"F9";
            when x"1EF" => DATA <= x"35";
            when x"1F0" => DATA <= x"8B";
            when x"1F1" => DATA <= x"80";
            when x"1F2" => DATA <= x"34";
            when x"1F3" => DATA <= x"01";
            when x"1F4" => DATA <= x"BD";
            when x"1F5" => DATA <= x"F9";
            when x"1F6" => DATA <= x"35";
            when x"1F7" => DATA <= x"1F";
            when x"1F8" => DATA <= x"89";
            when x"1F9" => DATA <= x"4F";
            when x"1FA" => DATA <= x"1F";
            when x"1FB" => DATA <= x"02";
            when x"1FC" => DATA <= x"BD";
            when x"1FD" => DATA <= x"F9";
            when x"1FE" => DATA <= x"35";
            when x"1FF" => DATA <= x"1E";
            when x"200" => DATA <= x"89";
            when x"201" => DATA <= x"1F";
            when x"202" => DATA <= x"01";
            when x"203" => DATA <= x"35";
            when x"204" => DATA <= x"87";
            when x"205" => DATA <= x"8E";
            when x"206" => DATA <= x"00";
            when x"207" => DATA <= x"00";
            when x"208" => DATA <= x"39";
            when x"209" => DATA <= x"BE";
            when x"20A" => DATA <= x"FF";
            when x"20B" => DATA <= x"88";
            when x"20C" => DATA <= x"39";
            when x"20D" => DATA <= x"BE";
            when x"20E" => DATA <= x"FF";
            when x"20F" => DATA <= x"8A";
            when x"210" => DATA <= x"39";
            when x"211" => DATA <= x"4D";
            when x"212" => DATA <= x"27";
            when x"213" => DATA <= x"60";
            when x"214" => DATA <= x"34";
            when x"215" => DATA <= x"26";
            when x"216" => DATA <= x"34";
            when x"217" => DATA <= x"10";
            when x"218" => DATA <= x"1F";
            when x"219" => DATA <= x"89";
            when x"21A" => DATA <= x"86";
            when x"21B" => DATA <= x"08";
            when x"21C" => DATA <= x"BD";
            when x"21D" => DATA <= x"FB";
            when x"21E" => DATA <= x"CA";
            when x"21F" => DATA <= x"1F";
            when x"220" => DATA <= x"98";
            when x"221" => DATA <= x"BD";
            when x"222" => DATA <= x"FB";
            when x"223" => DATA <= x"CA";
            when x"224" => DATA <= x"C1";
            when x"225" => DATA <= x"80";
            when x"226" => DATA <= x"24";
            when x"227" => DATA <= x"04";
            when x"228" => DATA <= x"A6";
            when x"229" => DATA <= x"84";
            when x"22A" => DATA <= x"20";
            when x"22B" => DATA <= x"0C";
            when x"22C" => DATA <= x"86";
            when x"22D" => DATA <= x"10";
            when x"22E" => DATA <= x"C1";
            when x"22F" => DATA <= x"15";
            when x"230" => DATA <= x"24";
            when x"231" => DATA <= x"06";
            when x"232" => DATA <= x"8E";
            when x"233" => DATA <= x"FA";
            when x"234" => DATA <= x"A5";
            when x"235" => DATA <= x"3A";
            when x"236" => DATA <= x"A6";
            when x"237" => DATA <= x"84";
            when x"238" => DATA <= x"35";
            when x"239" => DATA <= x"10";
            when x"23A" => DATA <= x"BD";
            when x"23B" => DATA <= x"FB";
            when x"23C" => DATA <= x"CA";
            when x"23D" => DATA <= x"1F";
            when x"23E" => DATA <= x"02";
            when x"23F" => DATA <= x"1E";
            when x"240" => DATA <= x"89";
            when x"241" => DATA <= x"4F";
            when x"242" => DATA <= x"1E";
            when x"243" => DATA <= x"02";
            when x"244" => DATA <= x"4A";
            when x"245" => DATA <= x"2B";
            when x"246" => DATA <= x"03";
            when x"247" => DATA <= x"BD";
            when x"248" => DATA <= x"FB";
            when x"249" => DATA <= x"98";
            when x"24A" => DATA <= x"34";
            when x"24B" => DATA <= x"10";
            when x"24C" => DATA <= x"C1";
            when x"24D" => DATA <= x"80";
            when x"24E" => DATA <= x"24";
            when x"24F" => DATA <= x"04";
            when x"250" => DATA <= x"A6";
            when x"251" => DATA <= x"01";
            when x"252" => DATA <= x"20";
            when x"253" => DATA <= x"0C";
            when x"254" => DATA <= x"86";
            when x"255" => DATA <= x"10";
            when x"256" => DATA <= x"C1";
            when x"257" => DATA <= x"15";
            when x"258" => DATA <= x"24";
            when x"259" => DATA <= x"06";
            when x"25A" => DATA <= x"8E";
            when x"25B" => DATA <= x"FA";
            when x"25C" => DATA <= x"B9";
            when x"25D" => DATA <= x"3A";
            when x"25E" => DATA <= x"A6";
            when x"25F" => DATA <= x"84";
            when x"260" => DATA <= x"35";
            when x"261" => DATA <= x"10";
            when x"262" => DATA <= x"BD";
            when x"263" => DATA <= x"FB";
            when x"264" => DATA <= x"CA";
            when x"265" => DATA <= x"1F";
            when x"266" => DATA <= x"02";
            when x"267" => DATA <= x"1E";
            when x"268" => DATA <= x"89";
            when x"269" => DATA <= x"4F";
            when x"26A" => DATA <= x"1E";
            when x"26B" => DATA <= x"02";
            when x"26C" => DATA <= x"4A";
            when x"26D" => DATA <= x"2B";
            when x"26E" => DATA <= x"03";
            when x"26F" => DATA <= x"BD";
            when x"270" => DATA <= x"FB";
            when x"271" => DATA <= x"A8";
            when x"272" => DATA <= x"35";
            when x"273" => DATA <= x"A6";
            when x"274" => DATA <= x"86";
            when x"275" => DATA <= x"0A";
            when x"276" => DATA <= x"BD";
            when x"277" => DATA <= x"FB";
            when x"278" => DATA <= x"CA";
            when x"279" => DATA <= x"30";
            when x"27A" => DATA <= x"02";
            when x"27B" => DATA <= x"10";
            when x"27C" => DATA <= x"8E";
            when x"27D" => DATA <= x"00";
            when x"27E" => DATA <= x"03";
            when x"27F" => DATA <= x"BD";
            when x"280" => DATA <= x"FB";
            when x"281" => DATA <= x"98";
            when x"282" => DATA <= x"30";
            when x"283" => DATA <= x"1E";
            when x"284" => DATA <= x"86";
            when x"285" => DATA <= x"07";
            when x"286" => DATA <= x"BD";
            when x"287" => DATA <= x"FB";
            when x"288" => DATA <= x"CA";
            when x"289" => DATA <= x"4F";
            when x"28A" => DATA <= x"BD";
            when x"28B" => DATA <= x"FB";
            when x"28C" => DATA <= x"CA";
            when x"28D" => DATA <= x"BD";
            when x"28E" => DATA <= x"F9";
            when x"28F" => DATA <= x"35";
            when x"290" => DATA <= x"8B";
            when x"291" => DATA <= x"80";
            when x"292" => DATA <= x"25";
            when x"293" => DATA <= x"11";
            when x"294" => DATA <= x"AE";
            when x"295" => DATA <= x"84";
            when x"296" => DATA <= x"BD";
            when x"297" => DATA <= x"F9";
            when x"298" => DATA <= x"35";
            when x"299" => DATA <= x"A7";
            when x"29A" => DATA <= x"80";
            when x"29B" => DATA <= x"31";
            when x"29C" => DATA <= x"21";
            when x"29D" => DATA <= x"81";
            when x"29E" => DATA <= x"0D";
            when x"29F" => DATA <= x"26";
            when x"2A0" => DATA <= x"F5";
            when x"2A1" => DATA <= x"31";
            when x"2A2" => DATA <= x"3F";
            when x"2A3" => DATA <= x"1C";
            when x"2A4" => DATA <= x"FE";
            when x"2A5" => DATA <= x"39";
            when x"2A6" => DATA <= x"00";
            when x"2A7" => DATA <= x"05";
            when x"2A8" => DATA <= x"00";
            when x"2A9" => DATA <= x"05";
            when x"2AA" => DATA <= x"04";
            when x"2AB" => DATA <= x"05";
            when x"2AC" => DATA <= x"08";
            when x"2AD" => DATA <= x"0E";
            when x"2AE" => DATA <= x"04";
            when x"2AF" => DATA <= x"01";
            when x"2B0" => DATA <= x"01";
            when x"2B1" => DATA <= x"05";
            when x"2B2" => DATA <= x"00";
            when x"2B3" => DATA <= x"01";
            when x"2B4" => DATA <= x"20";
            when x"2B5" => DATA <= x"10";
            when x"2B6" => DATA <= x"0D";
            when x"2B7" => DATA <= x"00";
            when x"2B8" => DATA <= x"04";
            when x"2B9" => DATA <= x"80";
            when x"2BA" => DATA <= x"05";
            when x"2BB" => DATA <= x"00";
            when x"2BC" => DATA <= x"05";
            when x"2BD" => DATA <= x"00";
            when x"2BE" => DATA <= x"05";
            when x"2BF" => DATA <= x"00";
            when x"2C0" => DATA <= x"00";
            when x"2C1" => DATA <= x"00";
            when x"2C2" => DATA <= x"05";
            when x"2C3" => DATA <= x"09";
            when x"2C4" => DATA <= x"05";
            when x"2C5" => DATA <= x"00";
            when x"2C6" => DATA <= x"08";
            when x"2C7" => DATA <= x"19";
            when x"2C8" => DATA <= x"00";
            when x"2C9" => DATA <= x"01";
            when x"2CA" => DATA <= x"0D";
            when x"2CB" => DATA <= x"80";
            when x"2CC" => DATA <= x"04";
            when x"2CD" => DATA <= x"80";
            when x"2CE" => DATA <= x"34";
            when x"2CF" => DATA <= x"26";
            when x"2D0" => DATA <= x"86";
            when x"2D1" => DATA <= x"0C";
            when x"2D2" => DATA <= x"BD";
            when x"2D3" => DATA <= x"FB";
            when x"2D4" => DATA <= x"CA";
            when x"2D5" => DATA <= x"1F";
            when x"2D6" => DATA <= x"20";
            when x"2D7" => DATA <= x"BD";
            when x"2D8" => DATA <= x"FB";
            when x"2D9" => DATA <= x"C8";
            when x"2DA" => DATA <= x"10";
            when x"2DB" => DATA <= x"8E";
            when x"2DC" => DATA <= x"00";
            when x"2DD" => DATA <= x"04";
            when x"2DE" => DATA <= x"BD";
            when x"2DF" => DATA <= x"FB";
            when x"2E0" => DATA <= x"98";
            when x"2E1" => DATA <= x"35";
            when x"2E2" => DATA <= x"06";
            when x"2E3" => DATA <= x"BD";
            when x"2E4" => DATA <= x"FB";
            when x"2E5" => DATA <= x"CA";
            when x"2E6" => DATA <= x"BD";
            when x"2E7" => DATA <= x"F9";
            when x"2E8" => DATA <= x"35";
            when x"2E9" => DATA <= x"34";
            when x"2EA" => DATA <= x"02";
            when x"2EB" => DATA <= x"10";
            when x"2EC" => DATA <= x"8E";
            when x"2ED" => DATA <= x"00";
            when x"2EE" => DATA <= x"04";
            when x"2EF" => DATA <= x"BD";
            when x"2F0" => DATA <= x"FB";
            when x"2F1" => DATA <= x"A8";
            when x"2F2" => DATA <= x"35";
            when x"2F3" => DATA <= x"A2";
            when x"2F4" => DATA <= x"86";
            when x"2F5" => DATA <= x"0E";
            when x"2F6" => DATA <= x"BD";
            when x"2F7" => DATA <= x"FB";
            when x"2F8" => DATA <= x"CA";
            when x"2F9" => DATA <= x"34";
            when x"2FA" => DATA <= x"06";
            when x"2FB" => DATA <= x"1F";
            when x"2FC" => DATA <= x"20";
            when x"2FD" => DATA <= x"BD";
            when x"2FE" => DATA <= x"FB";
            when x"2FF" => DATA <= x"C8";
            when x"300" => DATA <= x"35";
            when x"301" => DATA <= x"06";
            when x"302" => DATA <= x"7E";
            when x"303" => DATA <= x"F9";
            when x"304" => DATA <= x"31";
            when x"305" => DATA <= x"34";
            when x"306" => DATA <= x"06";
            when x"307" => DATA <= x"86";
            when x"308" => DATA <= x"10";
            when x"309" => DATA <= x"BD";
            when x"30A" => DATA <= x"FB";
            when x"30B" => DATA <= x"CA";
            when x"30C" => DATA <= x"1F";
            when x"30D" => DATA <= x"20";
            when x"30E" => DATA <= x"BD";
            when x"30F" => DATA <= x"FB";
            when x"310" => DATA <= x"C8";
            when x"311" => DATA <= x"35";
            when x"312" => DATA <= x"06";
            when x"313" => DATA <= x"34";
            when x"314" => DATA <= x"06";
            when x"315" => DATA <= x"BD";
            when x"316" => DATA <= x"FB";
            when x"317" => DATA <= x"CA";
            when x"318" => DATA <= x"BD";
            when x"319" => DATA <= x"F9";
            when x"31A" => DATA <= x"35";
            when x"31B" => DATA <= x"35";
            when x"31C" => DATA <= x"86";
            when x"31D" => DATA <= x"34";
            when x"31E" => DATA <= x"06";
            when x"31F" => DATA <= x"86";
            when x"320" => DATA <= x"12";
            when x"321" => DATA <= x"BD";
            when x"322" => DATA <= x"FB";
            when x"323" => DATA <= x"CA";
            when x"324" => DATA <= x"35";
            when x"325" => DATA <= x"06";
            when x"326" => DATA <= x"BD";
            when x"327" => DATA <= x"FB";
            when x"328" => DATA <= x"CA";
            when x"329" => DATA <= x"81";
            when x"32A" => DATA <= x"00";
            when x"32B" => DATA <= x"27";
            when x"32C" => DATA <= x"06";
            when x"32D" => DATA <= x"BD";
            when x"32E" => DATA <= x"FB";
            when x"32F" => DATA <= x"8F";
            when x"330" => DATA <= x"7E";
            when x"331" => DATA <= x"F9";
            when x"332" => DATA <= x"35";
            when x"333" => DATA <= x"34";
            when x"334" => DATA <= x"04";
            when x"335" => DATA <= x"1F";
            when x"336" => DATA <= x"20";
            when x"337" => DATA <= x"BD";
            when x"338" => DATA <= x"FB";
            when x"339" => DATA <= x"C8";
            when x"33A" => DATA <= x"BD";
            when x"33B" => DATA <= x"F9";
            when x"33C" => DATA <= x"35";
            when x"33D" => DATA <= x"4F";
            when x"33E" => DATA <= x"35";
            when x"33F" => DATA <= x"84";
            when x"340" => DATA <= x"34";
            when x"341" => DATA <= x"32";
            when x"342" => DATA <= x"86";
            when x"343" => DATA <= x"14";
            when x"344" => DATA <= x"BD";
            when x"345" => DATA <= x"FB";
            when x"346" => DATA <= x"CA";
            when x"347" => DATA <= x"30";
            when x"348" => DATA <= x"02";
            when x"349" => DATA <= x"10";
            when x"34A" => DATA <= x"8E";
            when x"34B" => DATA <= x"00";
            when x"34C" => DATA <= x"10";
            when x"34D" => DATA <= x"BD";
            when x"34E" => DATA <= x"FB";
            when x"34F" => DATA <= x"98";
            when x"350" => DATA <= x"30";
            when x"351" => DATA <= x"1E";
            when x"352" => DATA <= x"AE";
            when x"353" => DATA <= x"84";
            when x"354" => DATA <= x"BD";
            when x"355" => DATA <= x"FB";
            when x"356" => DATA <= x"8F";
            when x"357" => DATA <= x"35";
            when x"358" => DATA <= x"02";
            when x"359" => DATA <= x"BD";
            when x"35A" => DATA <= x"FB";
            when x"35B" => DATA <= x"CA";
            when x"35C" => DATA <= x"BD";
            when x"35D" => DATA <= x"F9";
            when x"35E" => DATA <= x"35";
            when x"35F" => DATA <= x"35";
            when x"360" => DATA <= x"10";
            when x"361" => DATA <= x"34";
            when x"362" => DATA <= x"02";
            when x"363" => DATA <= x"30";
            when x"364" => DATA <= x"02";
            when x"365" => DATA <= x"10";
            when x"366" => DATA <= x"8E";
            when x"367" => DATA <= x"00";
            when x"368" => DATA <= x"10";
            when x"369" => DATA <= x"BD";
            when x"36A" => DATA <= x"FB";
            when x"36B" => DATA <= x"A8";
            when x"36C" => DATA <= x"35";
            when x"36D" => DATA <= x"A2";
            when x"36E" => DATA <= x"34";
            when x"36F" => DATA <= x"20";
            when x"370" => DATA <= x"34";
            when x"371" => DATA <= x"02";
            when x"372" => DATA <= x"86";
            when x"373" => DATA <= x"16";
            when x"374" => DATA <= x"BD";
            when x"375" => DATA <= x"FB";
            when x"376" => DATA <= x"CA";
            when x"377" => DATA <= x"10";
            when x"378" => DATA <= x"8E";
            when x"379" => DATA <= x"00";
            when x"37A" => DATA <= x"0D";
            when x"37B" => DATA <= x"BD";
            when x"37C" => DATA <= x"FB";
            when x"37D" => DATA <= x"98";
            when x"37E" => DATA <= x"35";
            when x"37F" => DATA <= x"02";
            when x"380" => DATA <= x"BD";
            when x"381" => DATA <= x"FB";
            when x"382" => DATA <= x"CA";
            when x"383" => DATA <= x"10";
            when x"384" => DATA <= x"8E";
            when x"385" => DATA <= x"00";
            when x"386" => DATA <= x"0D";
            when x"387" => DATA <= x"BD";
            when x"388" => DATA <= x"FB";
            when x"389" => DATA <= x"A8";
            when x"38A" => DATA <= x"35";
            when x"38B" => DATA <= x"20";
            when x"38C" => DATA <= x"7E";
            when x"38D" => DATA <= x"F9";
            when x"38E" => DATA <= x"31";
            when x"38F" => DATA <= x"A6";
            when x"390" => DATA <= x"80";
            when x"391" => DATA <= x"8D";
            when x"392" => DATA <= x"37";
            when x"393" => DATA <= x"81";
            when x"394" => DATA <= x"0D";
            when x"395" => DATA <= x"26";
            when x"396" => DATA <= x"F8";
            when x"397" => DATA <= x"39";
            when x"398" => DATA <= x"34";
            when x"399" => DATA <= x"04";
            when x"39A" => DATA <= x"1F";
            when x"39B" => DATA <= x"20";
            when x"39C" => DATA <= x"3A";
            when x"39D" => DATA <= x"35";
            when x"39E" => DATA <= x"04";
            when x"39F" => DATA <= x"A6";
            when x"3A0" => DATA <= x"82";
            when x"3A1" => DATA <= x"8D";
            when x"3A2" => DATA <= x"27";
            when x"3A3" => DATA <= x"31";
            when x"3A4" => DATA <= x"3F";
            when x"3A5" => DATA <= x"26";
            when x"3A6" => DATA <= x"F8";
            when x"3A7" => DATA <= x"39";
            when x"3A8" => DATA <= x"34";
            when x"3A9" => DATA <= x"04";
            when x"3AA" => DATA <= x"1F";
            when x"3AB" => DATA <= x"20";
            when x"3AC" => DATA <= x"3A";
            when x"3AD" => DATA <= x"35";
            when x"3AE" => DATA <= x"04";
            when x"3AF" => DATA <= x"BD";
            when x"3B0" => DATA <= x"F9";
            when x"3B1" => DATA <= x"35";
            when x"3B2" => DATA <= x"A7";
            when x"3B3" => DATA <= x"82";
            when x"3B4" => DATA <= x"31";
            when x"3B5" => DATA <= x"3F";
            when x"3B6" => DATA <= x"26";
            when x"3B7" => DATA <= x"F7";
            when x"3B8" => DATA <= x"39";
            when x"3B9" => DATA <= x"34";
            when x"3BA" => DATA <= x"02";
            when x"3BB" => DATA <= x"B6";
            when x"3BC" => DATA <= x"FE";
            when x"3BD" => DATA <= x"E0";
            when x"3BE" => DATA <= x"84";
            when x"3BF" => DATA <= x"40";
            when x"3C0" => DATA <= x"27";
            when x"3C1" => DATA <= x"F9";
            when x"3C2" => DATA <= x"35";
            when x"3C3" => DATA <= x"02";
            when x"3C4" => DATA <= x"B7";
            when x"3C5" => DATA <= x"FE";
            when x"3C6" => DATA <= x"E1";
            when x"3C7" => DATA <= x"39";
            when x"3C8" => DATA <= x"1F";
            when x"3C9" => DATA <= x"98";
            when x"3CA" => DATA <= x"34";
            when x"3CB" => DATA <= x"02";
            when x"3CC" => DATA <= x"B6";
            when x"3CD" => DATA <= x"FE";
            when x"3CE" => DATA <= x"E2";
            when x"3CF" => DATA <= x"84";
            when x"3D0" => DATA <= x"40";
            when x"3D1" => DATA <= x"27";
            when x"3D2" => DATA <= x"F9";
            when x"3D3" => DATA <= x"35";
            when x"3D4" => DATA <= x"02";
            when x"3D5" => DATA <= x"B7";
            when x"3D6" => DATA <= x"FE";
            when x"3D7" => DATA <= x"E3";
            when x"3D8" => DATA <= x"39";
            when x"3D9" => DATA <= x"34";
            when x"3DA" => DATA <= x"02";
            when x"3DB" => DATA <= x"B6";
            when x"3DC" => DATA <= x"FE";
            when x"3DD" => DATA <= x"E6";
            when x"3DE" => DATA <= x"2B";
            when x"3DF" => DATA <= x"4F";
            when x"3E0" => DATA <= x"B6";
            when x"3E1" => DATA <= x"FE";
            when x"3E2" => DATA <= x"E0";
            when x"3E3" => DATA <= x"2B";
            when x"3E4" => DATA <= x"06";
            when x"3E5" => DATA <= x"35";
            when x"3E6" => DATA <= x"02";
            when x"3E7" => DATA <= x"6E";
            when x"3E8" => DATA <= x"9F";
            when x"3E9" => DATA <= x"FF";
            when x"3EA" => DATA <= x"B1";
            when x"3EB" => DATA <= x"B6";
            when x"3EC" => DATA <= x"FE";
            when x"3ED" => DATA <= x"E1";
            when x"3EE" => DATA <= x"2B";
            when x"3EF" => DATA <= x"1B";
            when x"3F0" => DATA <= x"34";
            when x"3F1" => DATA <= x"74";
            when x"3F2" => DATA <= x"8D";
            when x"3F3" => DATA <= x"1E";
            when x"3F4" => DATA <= x"1F";
            when x"3F5" => DATA <= x"89";
            when x"3F6" => DATA <= x"4F";
            when x"3F7" => DATA <= x"1F";
            when x"3F8" => DATA <= x"02";
            when x"3F9" => DATA <= x"8D";
            when x"3FA" => DATA <= x"17";
            when x"3FB" => DATA <= x"1F";
            when x"3FC" => DATA <= x"89";
            when x"3FD" => DATA <= x"4F";
            when x"3FE" => DATA <= x"1F";
            when x"3FF" => DATA <= x"01";
            when x"400" => DATA <= x"8D";
            when x"401" => DATA <= x"10";
            when x"402" => DATA <= x"AD";
            when x"403" => DATA <= x"9F";
            when x"404" => DATA <= x"FF";
            when x"405" => DATA <= x"FC";
            when x"406" => DATA <= x"35";
            when x"407" => DATA <= x"74";
            when x"408" => DATA <= x"35";
            when x"409" => DATA <= x"02";
            when x"40A" => DATA <= x"3B";
            when x"40B" => DATA <= x"49";
            when x"40C" => DATA <= x"B7";
            when x"40D" => DATA <= x"FF";
            when x"40E" => DATA <= x"80";
            when x"40F" => DATA <= x"35";
            when x"410" => DATA <= x"02";
            when x"411" => DATA <= x"3B";
            when x"412" => DATA <= x"B6";
            when x"413" => DATA <= x"FE";
            when x"414" => DATA <= x"E6";
            when x"415" => DATA <= x"2B";
            when x"416" => DATA <= x"02";
            when x"417" => DATA <= x"8D";
            when x"418" => DATA <= x"12";
            when x"419" => DATA <= x"B6";
            when x"41A" => DATA <= x"FE";
            when x"41B" => DATA <= x"E0";
            when x"41C" => DATA <= x"2A";
            when x"41D" => DATA <= x"F4";
            when x"41E" => DATA <= x"B6";
            when x"41F" => DATA <= x"FE";
            when x"420" => DATA <= x"E1";
            when x"421" => DATA <= x"39";
            when x"422" => DATA <= x"B6";
            when x"423" => DATA <= x"FE";
            when x"424" => DATA <= x"E6";
            when x"425" => DATA <= x"2A";
            when x"426" => DATA <= x"FB";
            when x"427" => DATA <= x"B6";
            when x"428" => DATA <= x"FE";
            when x"429" => DATA <= x"E7";
            when x"42A" => DATA <= x"39";
            when x"42B" => DATA <= x"1C";
            when x"42C" => DATA <= x"7F";
            when x"42D" => DATA <= x"34";
            when x"42E" => DATA <= x"01";
            when x"42F" => DATA <= x"B6";
            when x"430" => DATA <= x"FE";
            when x"431" => DATA <= x"E7";
            when x"432" => DATA <= x"2A";
            when x"433" => DATA <= x"20";
            when x"434" => DATA <= x"10";
            when x"435" => DATA <= x"CE";
            when x"436" => DATA <= x"FF";
            when x"437" => DATA <= x"80";
            when x"438" => DATA <= x"8E";
            when x"439" => DATA <= x"FF";
            when x"43A" => DATA <= x"00";
            when x"43B" => DATA <= x"BD";
            when x"43C" => DATA <= x"F9";
            when x"43D" => DATA <= x"35";
            when x"43E" => DATA <= x"86";
            when x"43F" => DATA <= x"3F";
            when x"440" => DATA <= x"A7";
            when x"441" => DATA <= x"80";
            when x"442" => DATA <= x"BD";
            when x"443" => DATA <= x"F9";
            when x"444" => DATA <= x"35";
            when x"445" => DATA <= x"A7";
            when x"446" => DATA <= x"80";
            when x"447" => DATA <= x"BD";
            when x"448" => DATA <= x"F9";
            when x"449" => DATA <= x"35";
            when x"44A" => DATA <= x"A7";
            when x"44B" => DATA <= x"80";
            when x"44C" => DATA <= x"26";
            when x"44D" => DATA <= x"F9";
            when x"44E" => DATA <= x"8E";
            when x"44F" => DATA <= x"FF";
            when x"450" => DATA <= x"01";
            when x"451" => DATA <= x"7E";
            when x"452" => DATA <= x"FF";
            when x"453" => DATA <= x"BC";
            when x"454" => DATA <= x"34";
            when x"455" => DATA <= x"02";
            when x"456" => DATA <= x"8D";
            when x"457" => DATA <= x"CA";
            when x"458" => DATA <= x"35";
            when x"459" => DATA <= x"02";
            when x"45A" => DATA <= x"81";
            when x"45B" => DATA <= x"05";
            when x"45C" => DATA <= x"26";
            when x"45D" => DATA <= x"06";
            when x"45E" => DATA <= x"7F";
            when x"45F" => DATA <= x"FF";
            when x"460" => DATA <= x"94";
            when x"461" => DATA <= x"35";
            when x"462" => DATA <= x"02";
            when x"463" => DATA <= x"3B";
            when x"464" => DATA <= x"34";
            when x"465" => DATA <= x"02";
            when x"466" => DATA <= x"8D";
            when x"467" => DATA <= x"BA";
            when x"468" => DATA <= x"B7";
            when x"469" => DATA <= x"FF";
            when x"46A" => DATA <= x"8C";
            when x"46B" => DATA <= x"8D";
            when x"46C" => DATA <= x"B5";
            when x"46D" => DATA <= x"B7";
            when x"46E" => DATA <= x"FF";
            when x"46F" => DATA <= x"8D";
            when x"470" => DATA <= x"8D";
            when x"471" => DATA <= x"B0";
            when x"472" => DATA <= x"B7";
            when x"473" => DATA <= x"FF";
            when x"474" => DATA <= x"8E";
            when x"475" => DATA <= x"8D";
            when x"476" => DATA <= x"AB";
            when x"477" => DATA <= x"B7";
            when x"478" => DATA <= x"FF";
            when x"479" => DATA <= x"8F";
            when x"47A" => DATA <= x"8D";
            when x"47B" => DATA <= x"A6";
            when x"47C" => DATA <= x"86";
            when x"47D" => DATA <= x"FF";
            when x"47E" => DATA <= x"B7";
            when x"47F" => DATA <= x"FF";
            when x"480" => DATA <= x"94";
            when x"481" => DATA <= x"1C";
            when x"482" => DATA <= x"BF";
            when x"483" => DATA <= x"A6";
            when x"484" => DATA <= x"E0";
            when x"485" => DATA <= x"27";
            when x"486" => DATA <= x"17";
            when x"487" => DATA <= x"81";
            when x"488" => DATA <= x"02";
            when x"489" => DATA <= x"25";
            when x"48A" => DATA <= x"27";
            when x"48B" => DATA <= x"27";
            when x"48C" => DATA <= x"39";
            when x"48D" => DATA <= x"81";
            when x"48E" => DATA <= x"04";
            when x"48F" => DATA <= x"25";
            when x"490" => DATA <= x"4C";
            when x"491" => DATA <= x"27";
            when x"492" => DATA <= x"61";
            when x"493" => DATA <= x"81";
            when x"494" => DATA <= x"07";
            when x"495" => DATA <= x"25";
            when x"496" => DATA <= x"66";
            when x"497" => DATA <= x"10";
            when x"498" => DATA <= x"27";
            when x"499" => DATA <= x"00";
            when x"49A" => DATA <= x"83";
            when x"49B" => DATA <= x"35";
            when x"49C" => DATA <= x"02";
            when x"49D" => DATA <= x"3B";
            when x"49E" => DATA <= x"BE";
            when x"49F" => DATA <= x"FF";
            when x"4A0" => DATA <= x"8E";
            when x"4A1" => DATA <= x"13";
            when x"4A2" => DATA <= x"A6";
            when x"4A3" => DATA <= x"80";
            when x"4A4" => DATA <= x"B7";
            when x"4A5" => DATA <= x"FE";
            when x"4A6" => DATA <= x"E5";
            when x"4A7" => DATA <= x"B6";
            when x"4A8" => DATA <= x"FF";
            when x"4A9" => DATA <= x"94";
            when x"4AA" => DATA <= x"26";
            when x"4AB" => DATA <= x"F5";
            when x"4AC" => DATA <= x"BF";
            when x"4AD" => DATA <= x"FF";
            when x"4AE" => DATA <= x"8E";
            when x"4AF" => DATA <= x"35";
            when x"4B0" => DATA <= x"02";
            when x"4B1" => DATA <= x"3B";
            when x"4B2" => DATA <= x"BE";
            when x"4B3" => DATA <= x"FF";
            when x"4B4" => DATA <= x"8E";
            when x"4B5" => DATA <= x"13";
            when x"4B6" => DATA <= x"B6";
            when x"4B7" => DATA <= x"FE";
            when x"4B8" => DATA <= x"E5";
            when x"4B9" => DATA <= x"A7";
            when x"4BA" => DATA <= x"80";
            when x"4BB" => DATA <= x"B6";
            when x"4BC" => DATA <= x"FF";
            when x"4BD" => DATA <= x"94";
            when x"4BE" => DATA <= x"26";
            when x"4BF" => DATA <= x"F5";
            when x"4C0" => DATA <= x"BF";
            when x"4C1" => DATA <= x"FF";
            when x"4C2" => DATA <= x"8E";
            when x"4C3" => DATA <= x"35";
            when x"4C4" => DATA <= x"02";
            when x"4C5" => DATA <= x"3B";
            when x"4C6" => DATA <= x"BE";
            when x"4C7" => DATA <= x"FF";
            when x"4C8" => DATA <= x"8E";
            when x"4C9" => DATA <= x"13";
            when x"4CA" => DATA <= x"EC";
            when x"4CB" => DATA <= x"81";
            when x"4CC" => DATA <= x"B7";
            when x"4CD" => DATA <= x"FE";
            when x"4CE" => DATA <= x"E5";
            when x"4CF" => DATA <= x"F7";
            when x"4D0" => DATA <= x"FE";
            when x"4D1" => DATA <= x"E5";
            when x"4D2" => DATA <= x"B6";
            when x"4D3" => DATA <= x"FF";
            when x"4D4" => DATA <= x"94";
            when x"4D5" => DATA <= x"26";
            when x"4D6" => DATA <= x"F2";
            when x"4D7" => DATA <= x"BF";
            when x"4D8" => DATA <= x"FF";
            when x"4D9" => DATA <= x"8E";
            when x"4DA" => DATA <= x"35";
            when x"4DB" => DATA <= x"02";
            when x"4DC" => DATA <= x"3B";
            when x"4DD" => DATA <= x"BE";
            when x"4DE" => DATA <= x"FF";
            when x"4DF" => DATA <= x"8E";
            when x"4E0" => DATA <= x"13";
            when x"4E1" => DATA <= x"B6";
            when x"4E2" => DATA <= x"FE";
            when x"4E3" => DATA <= x"E5";
            when x"4E4" => DATA <= x"F6";
            when x"4E5" => DATA <= x"FE";
            when x"4E6" => DATA <= x"E5";
            when x"4E7" => DATA <= x"ED";
            when x"4E8" => DATA <= x"81";
            when x"4E9" => DATA <= x"B6";
            when x"4EA" => DATA <= x"FF";
            when x"4EB" => DATA <= x"94";
            when x"4EC" => DATA <= x"26";
            when x"4ED" => DATA <= x"F2";
            when x"4EE" => DATA <= x"BF";
            when x"4EF" => DATA <= x"FF";
            when x"4F0" => DATA <= x"8E";
            when x"4F1" => DATA <= x"35";
            when x"4F2" => DATA <= x"02";
            when x"4F3" => DATA <= x"3B";
            when x"4F4" => DATA <= x"FC";
            when x"4F5" => DATA <= x"FF";
            when x"4F6" => DATA <= x"8E";
            when x"4F7" => DATA <= x"FD";
            when x"4F8" => DATA <= x"FF";
            when x"4F9" => DATA <= x"90";
            when x"4FA" => DATA <= x"35";
            when x"4FB" => DATA <= x"02";
            when x"4FC" => DATA <= x"3B";
            when x"4FD" => DATA <= x"34";
            when x"4FE" => DATA <= x"04";
            when x"4FF" => DATA <= x"BE";
            when x"500" => DATA <= x"FF";
            when x"501" => DATA <= x"8E";
            when x"502" => DATA <= x"5F";
            when x"503" => DATA <= x"B6";
            when x"504" => DATA <= x"FE";
            when x"505" => DATA <= x"E4";
            when x"506" => DATA <= x"84";
            when x"507" => DATA <= x"40";
            when x"508" => DATA <= x"27";
            when x"509" => DATA <= x"F9";
            when x"50A" => DATA <= x"B6";
            when x"50B" => DATA <= x"FE";
            when x"50C" => DATA <= x"E5";
            when x"50D" => DATA <= x"A7";
            when x"50E" => DATA <= x"85";
            when x"50F" => DATA <= x"5C";
            when x"510" => DATA <= x"26";
            when x"511" => DATA <= x"F1";
            when x"512" => DATA <= x"30";
            when x"513" => DATA <= x"89";
            when x"514" => DATA <= x"01";
            when x"515" => DATA <= x"00";
            when x"516" => DATA <= x"BF";
            when x"517" => DATA <= x"FF";
            when x"518" => DATA <= x"8E";
            when x"519" => DATA <= x"35";
            when x"51A" => DATA <= x"04";
            when x"51B" => DATA <= x"35";
            when x"51C" => DATA <= x"02";
            when x"51D" => DATA <= x"3B";
            when x"51E" => DATA <= x"34";
            when x"51F" => DATA <= x"04";
            when x"520" => DATA <= x"BE";
            when x"521" => DATA <= x"FF";
            when x"522" => DATA <= x"8E";
            when x"523" => DATA <= x"5F";
            when x"524" => DATA <= x"B6";
            when x"525" => DATA <= x"FE";
            when x"526" => DATA <= x"E4";
            when x"527" => DATA <= x"2A";
            when x"528" => DATA <= x"FB";
            when x"529" => DATA <= x"A6";
            when x"52A" => DATA <= x"85";
            when x"52B" => DATA <= x"B7";
            when x"52C" => DATA <= x"FE";
            when x"52D" => DATA <= x"E5";
            when x"52E" => DATA <= x"5C";
            when x"52F" => DATA <= x"26";
            when x"530" => DATA <= x"F3";
            when x"531" => DATA <= x"30";
            when x"532" => DATA <= x"89";
            when x"533" => DATA <= x"01";
            when x"534" => DATA <= x"00";
            when x"535" => DATA <= x"BF";
            when x"536" => DATA <= x"FF";
            when x"537" => DATA <= x"8E";
            when x"538" => DATA <= x"35";
            when x"539" => DATA <= x"04";
            when x"53A" => DATA <= x"35";
            when x"53B" => DATA <= x"02";
            when x"53C" => DATA <= x"3B";
            when x"53D" => DATA <= x"AE";
            when x"53E" => DATA <= x"6A";
            when x"53F" => DATA <= x"1C";
            when x"540" => DATA <= x"00";
            when x"541" => DATA <= x"BF";
            when x"542" => DATA <= x"FF";
            when x"543" => DATA <= x"82";
            when x"544" => DATA <= x"6E";
            when x"545" => DATA <= x"9F";
            when x"546" => DATA <= x"FF";
            when x"547" => DATA <= x"FA";
            when x"548" => DATA <= x"FF";
            when x"549" => DATA <= x"FF";
            when x"54A" => DATA <= x"FF";
            when x"54B" => DATA <= x"FF";
            when x"54C" => DATA <= x"FF";
            when x"54D" => DATA <= x"FF";
            when x"54E" => DATA <= x"FF";
            when x"54F" => DATA <= x"FF";
            when x"550" => DATA <= x"FF";
            when x"551" => DATA <= x"FF";
            when x"552" => DATA <= x"FF";
            when x"553" => DATA <= x"FF";
            when x"554" => DATA <= x"FF";
            when x"555" => DATA <= x"FF";
            when x"556" => DATA <= x"FF";
            when x"557" => DATA <= x"FF";
            when x"558" => DATA <= x"FF";
            when x"559" => DATA <= x"FF";
            when x"55A" => DATA <= x"FF";
            when x"55B" => DATA <= x"FF";
            when x"55C" => DATA <= x"FF";
            when x"55D" => DATA <= x"FF";
            when x"55E" => DATA <= x"FF";
            when x"55F" => DATA <= x"FF";
            when x"560" => DATA <= x"FF";
            when x"561" => DATA <= x"FF";
            when x"562" => DATA <= x"FF";
            when x"563" => DATA <= x"FF";
            when x"564" => DATA <= x"FF";
            when x"565" => DATA <= x"FF";
            when x"566" => DATA <= x"FF";
            when x"567" => DATA <= x"FF";
            when x"568" => DATA <= x"FF";
            when x"569" => DATA <= x"FF";
            when x"56A" => DATA <= x"FF";
            when x"56B" => DATA <= x"FF";
            when x"56C" => DATA <= x"FF";
            when x"56D" => DATA <= x"FF";
            when x"56E" => DATA <= x"FF";
            when x"56F" => DATA <= x"FF";
            when x"570" => DATA <= x"FF";
            when x"571" => DATA <= x"FF";
            when x"572" => DATA <= x"FF";
            when x"573" => DATA <= x"FF";
            when x"574" => DATA <= x"FF";
            when x"575" => DATA <= x"FF";
            when x"576" => DATA <= x"FF";
            when x"577" => DATA <= x"FF";
            when x"578" => DATA <= x"FF";
            when x"579" => DATA <= x"FF";
            when x"57A" => DATA <= x"FF";
            when x"57B" => DATA <= x"FF";
            when x"57C" => DATA <= x"FF";
            when x"57D" => DATA <= x"FF";
            when x"57E" => DATA <= x"FF";
            when x"57F" => DATA <= x"FF";
            when x"580" => DATA <= x"FF";
            when x"581" => DATA <= x"FF";
            when x"582" => DATA <= x"FF";
            when x"583" => DATA <= x"FF";
            when x"584" => DATA <= x"FF";
            when x"585" => DATA <= x"FF";
            when x"586" => DATA <= x"FF";
            when x"587" => DATA <= x"FF";
            when x"588" => DATA <= x"FF";
            when x"589" => DATA <= x"FF";
            when x"58A" => DATA <= x"FF";
            when x"58B" => DATA <= x"FF";
            when x"58C" => DATA <= x"FF";
            when x"58D" => DATA <= x"FF";
            when x"58E" => DATA <= x"FF";
            when x"58F" => DATA <= x"FF";
            when x"590" => DATA <= x"FF";
            when x"591" => DATA <= x"FF";
            when x"592" => DATA <= x"FF";
            when x"593" => DATA <= x"FF";
            when x"594" => DATA <= x"FF";
            when x"595" => DATA <= x"FF";
            when x"596" => DATA <= x"FF";
            when x"597" => DATA <= x"FF";
            when x"598" => DATA <= x"FF";
            when x"599" => DATA <= x"FF";
            when x"59A" => DATA <= x"FF";
            when x"59B" => DATA <= x"FF";
            when x"59C" => DATA <= x"FF";
            when x"59D" => DATA <= x"FF";
            when x"59E" => DATA <= x"FF";
            when x"59F" => DATA <= x"FF";
            when x"5A0" => DATA <= x"FF";
            when x"5A1" => DATA <= x"FF";
            when x"5A2" => DATA <= x"FF";
            when x"5A3" => DATA <= x"FF";
            when x"5A4" => DATA <= x"FF";
            when x"5A5" => DATA <= x"FF";
            when x"5A6" => DATA <= x"FF";
            when x"5A7" => DATA <= x"FF";
            when x"5A8" => DATA <= x"FF";
            when x"5A9" => DATA <= x"FF";
            when x"5AA" => DATA <= x"FF";
            when x"5AB" => DATA <= x"FF";
            when x"5AC" => DATA <= x"FF";
            when x"5AD" => DATA <= x"FF";
            when x"5AE" => DATA <= x"FF";
            when x"5AF" => DATA <= x"FF";
            when x"5B0" => DATA <= x"FF";
            when x"5B1" => DATA <= x"FF";
            when x"5B2" => DATA <= x"FF";
            when x"5B3" => DATA <= x"FF";
            when x"5B4" => DATA <= x"FF";
            when x"5B5" => DATA <= x"FF";
            when x"5B6" => DATA <= x"FF";
            when x"5B7" => DATA <= x"FF";
            when x"5B8" => DATA <= x"FF";
            when x"5B9" => DATA <= x"FF";
            when x"5BA" => DATA <= x"FF";
            when x"5BB" => DATA <= x"FF";
            when x"5BC" => DATA <= x"FF";
            when x"5BD" => DATA <= x"FF";
            when x"5BE" => DATA <= x"FF";
            when x"5BF" => DATA <= x"FF";
            when x"5C0" => DATA <= x"FF";
            when x"5C1" => DATA <= x"FF";
            when x"5C2" => DATA <= x"FF";
            when x"5C3" => DATA <= x"FF";
            when x"5C4" => DATA <= x"FF";
            when x"5C5" => DATA <= x"FF";
            when x"5C6" => DATA <= x"FF";
            when x"5C7" => DATA <= x"FF";
            when x"5C8" => DATA <= x"FF";
            when x"5C9" => DATA <= x"FF";
            when x"5CA" => DATA <= x"FF";
            when x"5CB" => DATA <= x"FF";
            when x"5CC" => DATA <= x"FF";
            when x"5CD" => DATA <= x"FF";
            when x"5CE" => DATA <= x"FF";
            when x"5CF" => DATA <= x"FF";
            when x"5D0" => DATA <= x"FF";
            when x"5D1" => DATA <= x"FF";
            when x"5D2" => DATA <= x"FF";
            when x"5D3" => DATA <= x"FF";
            when x"5D4" => DATA <= x"FF";
            when x"5D5" => DATA <= x"FF";
            when x"5D6" => DATA <= x"FF";
            when x"5D7" => DATA <= x"FF";
            when x"5D8" => DATA <= x"FF";
            when x"5D9" => DATA <= x"FF";
            when x"5DA" => DATA <= x"FF";
            when x"5DB" => DATA <= x"FF";
            when x"5DC" => DATA <= x"FF";
            when x"5DD" => DATA <= x"FF";
            when x"5DE" => DATA <= x"FF";
            when x"5DF" => DATA <= x"FF";
            when x"5E0" => DATA <= x"FF";
            when x"5E1" => DATA <= x"FF";
            when x"5E2" => DATA <= x"FF";
            when x"5E3" => DATA <= x"FF";
            when x"5E4" => DATA <= x"FF";
            when x"5E5" => DATA <= x"FF";
            when x"5E6" => DATA <= x"FF";
            when x"5E7" => DATA <= x"FF";
            when x"5E8" => DATA <= x"FF";
            when x"5E9" => DATA <= x"FF";
            when x"5EA" => DATA <= x"FF";
            when x"5EB" => DATA <= x"FF";
            when x"5EC" => DATA <= x"FF";
            when x"5ED" => DATA <= x"FF";
            when x"5EE" => DATA <= x"FF";
            when x"5EF" => DATA <= x"FF";
            when x"5F0" => DATA <= x"FF";
            when x"5F1" => DATA <= x"FF";
            when x"5F2" => DATA <= x"FF";
            when x"5F3" => DATA <= x"FF";
            when x"5F4" => DATA <= x"FF";
            when x"5F5" => DATA <= x"FF";
            when x"5F6" => DATA <= x"FF";
            when x"5F7" => DATA <= x"FF";
            when x"5F8" => DATA <= x"FF";
            when x"5F9" => DATA <= x"FF";
            when x"5FA" => DATA <= x"FF";
            when x"5FB" => DATA <= x"FF";
            when x"5FC" => DATA <= x"FF";
            when x"5FD" => DATA <= x"FF";
            when x"5FE" => DATA <= x"FF";
            when x"5FF" => DATA <= x"FF";
            when x"600" => DATA <= x"FF";
            when x"601" => DATA <= x"FF";
            when x"602" => DATA <= x"FF";
            when x"603" => DATA <= x"FF";
            when x"604" => DATA <= x"FF";
            when x"605" => DATA <= x"FF";
            when x"606" => DATA <= x"FF";
            when x"607" => DATA <= x"FF";
            when x"608" => DATA <= x"FF";
            when x"609" => DATA <= x"FF";
            when x"60A" => DATA <= x"FF";
            when x"60B" => DATA <= x"FF";
            when x"60C" => DATA <= x"FF";
            when x"60D" => DATA <= x"FF";
            when x"60E" => DATA <= x"FF";
            when x"60F" => DATA <= x"FF";
            when x"610" => DATA <= x"FF";
            when x"611" => DATA <= x"FF";
            when x"612" => DATA <= x"FF";
            when x"613" => DATA <= x"FF";
            when x"614" => DATA <= x"FF";
            when x"615" => DATA <= x"FF";
            when x"616" => DATA <= x"FF";
            when x"617" => DATA <= x"FF";
            when x"618" => DATA <= x"FF";
            when x"619" => DATA <= x"FF";
            when x"61A" => DATA <= x"FF";
            when x"61B" => DATA <= x"FF";
            when x"61C" => DATA <= x"FF";
            when x"61D" => DATA <= x"FF";
            when x"61E" => DATA <= x"FF";
            when x"61F" => DATA <= x"FF";
            when x"620" => DATA <= x"FF";
            when x"621" => DATA <= x"FF";
            when x"622" => DATA <= x"FF";
            when x"623" => DATA <= x"FF";
            when x"624" => DATA <= x"FF";
            when x"625" => DATA <= x"FF";
            when x"626" => DATA <= x"FF";
            when x"627" => DATA <= x"FF";
            when x"628" => DATA <= x"FF";
            when x"629" => DATA <= x"FF";
            when x"62A" => DATA <= x"FF";
            when x"62B" => DATA <= x"FF";
            when x"62C" => DATA <= x"FF";
            when x"62D" => DATA <= x"FF";
            when x"62E" => DATA <= x"FF";
            when x"62F" => DATA <= x"FF";
            when x"630" => DATA <= x"FF";
            when x"631" => DATA <= x"FF";
            when x"632" => DATA <= x"FF";
            when x"633" => DATA <= x"FF";
            when x"634" => DATA <= x"FF";
            when x"635" => DATA <= x"FF";
            when x"636" => DATA <= x"FF";
            when x"637" => DATA <= x"FF";
            when x"638" => DATA <= x"FF";
            when x"639" => DATA <= x"FF";
            when x"63A" => DATA <= x"FF";
            when x"63B" => DATA <= x"FF";
            when x"63C" => DATA <= x"FF";
            when x"63D" => DATA <= x"FF";
            when x"63E" => DATA <= x"FF";
            when x"63F" => DATA <= x"FF";
            when x"640" => DATA <= x"FF";
            when x"641" => DATA <= x"FF";
            when x"642" => DATA <= x"FF";
            when x"643" => DATA <= x"FF";
            when x"644" => DATA <= x"FF";
            when x"645" => DATA <= x"FF";
            when x"646" => DATA <= x"FF";
            when x"647" => DATA <= x"FF";
            when x"648" => DATA <= x"FF";
            when x"649" => DATA <= x"FF";
            when x"64A" => DATA <= x"FF";
            when x"64B" => DATA <= x"FF";
            when x"64C" => DATA <= x"FF";
            when x"64D" => DATA <= x"FF";
            when x"64E" => DATA <= x"FF";
            when x"64F" => DATA <= x"FF";
            when x"650" => DATA <= x"FF";
            when x"651" => DATA <= x"FF";
            when x"652" => DATA <= x"FF";
            when x"653" => DATA <= x"FF";
            when x"654" => DATA <= x"FF";
            when x"655" => DATA <= x"FF";
            when x"656" => DATA <= x"FF";
            when x"657" => DATA <= x"FF";
            when x"658" => DATA <= x"FF";
            when x"659" => DATA <= x"FF";
            when x"65A" => DATA <= x"FF";
            when x"65B" => DATA <= x"FF";
            when x"65C" => DATA <= x"FF";
            when x"65D" => DATA <= x"FF";
            when x"65E" => DATA <= x"FF";
            when x"65F" => DATA <= x"FF";
            when x"660" => DATA <= x"FF";
            when x"661" => DATA <= x"FF";
            when x"662" => DATA <= x"FF";
            when x"663" => DATA <= x"FF";
            when x"664" => DATA <= x"FF";
            when x"665" => DATA <= x"FF";
            when x"666" => DATA <= x"FF";
            when x"667" => DATA <= x"FF";
            when x"668" => DATA <= x"FF";
            when x"669" => DATA <= x"FF";
            when x"66A" => DATA <= x"FF";
            when x"66B" => DATA <= x"FF";
            when x"66C" => DATA <= x"FF";
            when x"66D" => DATA <= x"FF";
            when x"66E" => DATA <= x"FF";
            when x"66F" => DATA <= x"FF";
            when x"670" => DATA <= x"FF";
            when x"671" => DATA <= x"FF";
            when x"672" => DATA <= x"FF";
            when x"673" => DATA <= x"FF";
            when x"674" => DATA <= x"FF";
            when x"675" => DATA <= x"FF";
            when x"676" => DATA <= x"FF";
            when x"677" => DATA <= x"FF";
            when x"678" => DATA <= x"FF";
            when x"679" => DATA <= x"FF";
            when x"67A" => DATA <= x"FF";
            when x"67B" => DATA <= x"FF";
            when x"67C" => DATA <= x"FF";
            when x"67D" => DATA <= x"FF";
            when x"67E" => DATA <= x"FF";
            when x"67F" => DATA <= x"FF";
            when x"680" => DATA <= x"FF";
            when x"681" => DATA <= x"FF";
            when x"682" => DATA <= x"FF";
            when x"683" => DATA <= x"FF";
            when x"684" => DATA <= x"FF";
            when x"685" => DATA <= x"FF";
            when x"686" => DATA <= x"FF";
            when x"687" => DATA <= x"FF";
            when x"688" => DATA <= x"FF";
            when x"689" => DATA <= x"FF";
            when x"68A" => DATA <= x"FF";
            when x"68B" => DATA <= x"FF";
            when x"68C" => DATA <= x"FF";
            when x"68D" => DATA <= x"FF";
            when x"68E" => DATA <= x"FF";
            when x"68F" => DATA <= x"FF";
            when x"690" => DATA <= x"FF";
            when x"691" => DATA <= x"FF";
            when x"692" => DATA <= x"FF";
            when x"693" => DATA <= x"FF";
            when x"694" => DATA <= x"FF";
            when x"695" => DATA <= x"FF";
            when x"696" => DATA <= x"FF";
            when x"697" => DATA <= x"FF";
            when x"698" => DATA <= x"FF";
            when x"699" => DATA <= x"FF";
            when x"69A" => DATA <= x"FF";
            when x"69B" => DATA <= x"FF";
            when x"69C" => DATA <= x"FF";
            when x"69D" => DATA <= x"FF";
            when x"69E" => DATA <= x"FF";
            when x"69F" => DATA <= x"FF";
            when x"6A0" => DATA <= x"FF";
            when x"6A1" => DATA <= x"FF";
            when x"6A2" => DATA <= x"FF";
            when x"6A3" => DATA <= x"FF";
            when x"6A4" => DATA <= x"FF";
            when x"6A5" => DATA <= x"FF";
            when x"6A6" => DATA <= x"FF";
            when x"6A7" => DATA <= x"FF";
            when x"6A8" => DATA <= x"FF";
            when x"6A9" => DATA <= x"FF";
            when x"6AA" => DATA <= x"FF";
            when x"6AB" => DATA <= x"FF";
            when x"6AC" => DATA <= x"FF";
            when x"6AD" => DATA <= x"FF";
            when x"6AE" => DATA <= x"FF";
            when x"6AF" => DATA <= x"FF";
            when x"6B0" => DATA <= x"FF";
            when x"6B1" => DATA <= x"FF";
            when x"6B2" => DATA <= x"FF";
            when x"6B3" => DATA <= x"FF";
            when x"6B4" => DATA <= x"FF";
            when x"6B5" => DATA <= x"FF";
            when x"6B6" => DATA <= x"FF";
            when x"6B7" => DATA <= x"FF";
            when x"6B8" => DATA <= x"FF";
            when x"6B9" => DATA <= x"FF";
            when x"6BA" => DATA <= x"FF";
            when x"6BB" => DATA <= x"FF";
            when x"6BC" => DATA <= x"FF";
            when x"6BD" => DATA <= x"FF";
            when x"6BE" => DATA <= x"FF";
            when x"6BF" => DATA <= x"FF";
            when x"6C0" => DATA <= x"FF";
            when x"6C1" => DATA <= x"FF";
            when x"6C2" => DATA <= x"FF";
            when x"6C3" => DATA <= x"FF";
            when x"6C4" => DATA <= x"FF";
            when x"6C5" => DATA <= x"FF";
            when x"6C6" => DATA <= x"FF";
            when x"6C7" => DATA <= x"FF";
            when x"6C8" => DATA <= x"FF";
            when x"6C9" => DATA <= x"FF";
            when x"6CA" => DATA <= x"FF";
            when x"6CB" => DATA <= x"FF";
            when x"6CC" => DATA <= x"FF";
            when x"6CD" => DATA <= x"FF";
            when x"6CE" => DATA <= x"FF";
            when x"6CF" => DATA <= x"FF";
            when x"6D0" => DATA <= x"FF";
            when x"6D1" => DATA <= x"FF";
            when x"6D2" => DATA <= x"FF";
            when x"6D3" => DATA <= x"FF";
            when x"6D4" => DATA <= x"FF";
            when x"6D5" => DATA <= x"FF";
            when x"6D6" => DATA <= x"FF";
            when x"6D7" => DATA <= x"FF";
            when x"6D8" => DATA <= x"FF";
            when x"6D9" => DATA <= x"FF";
            when x"6DA" => DATA <= x"FF";
            when x"6DB" => DATA <= x"FF";
            when x"6DC" => DATA <= x"FF";
            when x"6DD" => DATA <= x"FF";
            when x"6DE" => DATA <= x"FF";
            when x"6DF" => DATA <= x"FF";
            when x"6E0" => DATA <= x"00";
            when x"6E1" => DATA <= x"00";
            when x"6E2" => DATA <= x"00";
            when x"6E3" => DATA <= x"00";
            when x"6E4" => DATA <= x"00";
            when x"6E5" => DATA <= x"00";
            when x"6E6" => DATA <= x"00";
            when x"6E7" => DATA <= x"00";
            when x"6E8" => DATA <= x"FF";
            when x"6E9" => DATA <= x"FF";
            when x"6EA" => DATA <= x"FF";
            when x"6EB" => DATA <= x"FF";
            when x"6EC" => DATA <= x"FF";
            when x"6ED" => DATA <= x"FF";
            when x"6EE" => DATA <= x"FF";
            when x"6EF" => DATA <= x"FF";
            when x"6F0" => DATA <= x"FD";
            when x"6F1" => DATA <= x"3C";
            when x"6F2" => DATA <= x"FD";
            when x"6F3" => DATA <= x"3C";
            when x"6F4" => DATA <= x"FD";
            when x"6F5" => DATA <= x"3C";
            when x"6F6" => DATA <= x"FB";
            when x"6F7" => DATA <= x"D9";
            when x"6F8" => DATA <= x"FD";
            when x"6F9" => DATA <= x"3C";
            when x"6FA" => DATA <= x"FD";
            when x"6FB" => DATA <= x"3D";
            when x"6FC" => DATA <= x"FD";
            when x"6FD" => DATA <= x"3C";
            when x"6FE" => DATA <= x"F8";
            when x"6FF" => DATA <= x"2D";
            when x"700" => DATA <= x"00";
            when x"701" => DATA <= x"00";
            when x"702" => DATA <= x"00";
            when x"703" => DATA <= x"00";
            when x"704" => DATA <= x"00";
            when x"705" => DATA <= x"00";
            when x"706" => DATA <= x"00";
            when x"707" => DATA <= x"00";
            when x"708" => DATA <= x"00";
            when x"709" => DATA <= x"00";
            when x"70A" => DATA <= x"00";
            when x"70B" => DATA <= x"00";
            when x"70C" => DATA <= x"00";
            when x"70D" => DATA <= x"00";
            when x"70E" => DATA <= x"00";
            when x"70F" => DATA <= x"00";
            when x"710" => DATA <= x"00";
            when x"711" => DATA <= x"00";
            when x"712" => DATA <= x"00";
            when x"713" => DATA <= x"00";
            when x"714" => DATA <= x"00";
            when x"715" => DATA <= x"00";
            when x"716" => DATA <= x"00";
            when x"717" => DATA <= x"00";
            when x"718" => DATA <= x"00";
            when x"719" => DATA <= x"00";
            when x"71A" => DATA <= x"00";
            when x"71B" => DATA <= x"00";
            when x"71C" => DATA <= x"00";
            when x"71D" => DATA <= x"00";
            when x"71E" => DATA <= x"00";
            when x"71F" => DATA <= x"00";
            when x"720" => DATA <= x"00";
            when x"721" => DATA <= x"00";
            when x"722" => DATA <= x"00";
            when x"723" => DATA <= x"00";
            when x"724" => DATA <= x"00";
            when x"725" => DATA <= x"00";
            when x"726" => DATA <= x"00";
            when x"727" => DATA <= x"00";
            when x"728" => DATA <= x"00";
            when x"729" => DATA <= x"00";
            when x"72A" => DATA <= x"00";
            when x"72B" => DATA <= x"00";
            when x"72C" => DATA <= x"00";
            when x"72D" => DATA <= x"00";
            when x"72E" => DATA <= x"00";
            when x"72F" => DATA <= x"00";
            when x"730" => DATA <= x"00";
            when x"731" => DATA <= x"00";
            when x"732" => DATA <= x"00";
            when x"733" => DATA <= x"00";
            when x"734" => DATA <= x"00";
            when x"735" => DATA <= x"00";
            when x"736" => DATA <= x"00";
            when x"737" => DATA <= x"00";
            when x"738" => DATA <= x"00";
            when x"739" => DATA <= x"00";
            when x"73A" => DATA <= x"00";
            when x"73B" => DATA <= x"00";
            when x"73C" => DATA <= x"00";
            when x"73D" => DATA <= x"00";
            when x"73E" => DATA <= x"00";
            when x"73F" => DATA <= x"00";
            when x"740" => DATA <= x"00";
            when x"741" => DATA <= x"00";
            when x"742" => DATA <= x"00";
            when x"743" => DATA <= x"00";
            when x"744" => DATA <= x"00";
            when x"745" => DATA <= x"00";
            when x"746" => DATA <= x"00";
            when x"747" => DATA <= x"00";
            when x"748" => DATA <= x"00";
            when x"749" => DATA <= x"00";
            when x"74A" => DATA <= x"00";
            when x"74B" => DATA <= x"00";
            when x"74C" => DATA <= x"00";
            when x"74D" => DATA <= x"00";
            when x"74E" => DATA <= x"00";
            when x"74F" => DATA <= x"00";
            when x"750" => DATA <= x"00";
            when x"751" => DATA <= x"00";
            when x"752" => DATA <= x"00";
            when x"753" => DATA <= x"00";
            when x"754" => DATA <= x"00";
            when x"755" => DATA <= x"00";
            when x"756" => DATA <= x"00";
            when x"757" => DATA <= x"00";
            when x"758" => DATA <= x"00";
            when x"759" => DATA <= x"00";
            when x"75A" => DATA <= x"00";
            when x"75B" => DATA <= x"00";
            when x"75C" => DATA <= x"00";
            when x"75D" => DATA <= x"00";
            when x"75E" => DATA <= x"00";
            when x"75F" => DATA <= x"00";
            when x"760" => DATA <= x"00";
            when x"761" => DATA <= x"00";
            when x"762" => DATA <= x"00";
            when x"763" => DATA <= x"00";
            when x"764" => DATA <= x"00";
            when x"765" => DATA <= x"00";
            when x"766" => DATA <= x"00";
            when x"767" => DATA <= x"00";
            when x"768" => DATA <= x"00";
            when x"769" => DATA <= x"00";
            when x"76A" => DATA <= x"00";
            when x"76B" => DATA <= x"00";
            when x"76C" => DATA <= x"00";
            when x"76D" => DATA <= x"00";
            when x"76E" => DATA <= x"00";
            when x"76F" => DATA <= x"00";
            when x"770" => DATA <= x"00";
            when x"771" => DATA <= x"00";
            when x"772" => DATA <= x"00";
            when x"773" => DATA <= x"00";
            when x"774" => DATA <= x"00";
            when x"775" => DATA <= x"00";
            when x"776" => DATA <= x"00";
            when x"777" => DATA <= x"00";
            when x"778" => DATA <= x"00";
            when x"779" => DATA <= x"00";
            when x"77A" => DATA <= x"00";
            when x"77B" => DATA <= x"00";
            when x"77C" => DATA <= x"00";
            when x"77D" => DATA <= x"00";
            when x"77E" => DATA <= x"00";
            when x"77F" => DATA <= x"00";
            when x"780" => DATA <= x"00";
            when x"781" => DATA <= x"00";
            when x"782" => DATA <= x"F8";
            when x"783" => DATA <= x"16";
            when x"784" => DATA <= x"F8";
            when x"785" => DATA <= x"A7";
            when x"786" => DATA <= x"F8";
            when x"787" => DATA <= x"16";
            when x"788" => DATA <= x"00";
            when x"789" => DATA <= x"00";
            when x"78A" => DATA <= x"F8";
            when x"78B" => DATA <= x"00";
            when x"78C" => DATA <= x"00";
            when x"78D" => DATA <= x"00";
            when x"78E" => DATA <= x"00";
            when x"78F" => DATA <= x"00";
            when x"790" => DATA <= x"F8";
            when x"791" => DATA <= x"00";
            when x"792" => DATA <= x"00";
            when x"793" => DATA <= x"00";
            when x"794" => DATA <= x"00";
            when x"795" => DATA <= x"7E";
            when x"796" => DATA <= x"F9";
            when x"797" => DATA <= x"4D";
            when x"798" => DATA <= x"7E";
            when x"799" => DATA <= x"F9";
            when x"79A" => DATA <= x"4D";
            when x"79B" => DATA <= x"7E";
            when x"79C" => DATA <= x"F9";
            when x"79D" => DATA <= x"4D";
            when x"79E" => DATA <= x"7E";
            when x"79F" => DATA <= x"F9";
            when x"7A0" => DATA <= x"4D";
            when x"7A1" => DATA <= x"7E";
            when x"7A2" => DATA <= x"F9";
            when x"7A3" => DATA <= x"4D";
            when x"7A4" => DATA <= x"7E";
            when x"7A5" => DATA <= x"F9";
            when x"7A6" => DATA <= x"4D";
            when x"7A7" => DATA <= x"7E";
            when x"7A8" => DATA <= x"F8";
            when x"7A9" => DATA <= x"67";
            when x"7AA" => DATA <= x"7E";
            when x"7AB" => DATA <= x"F9";
            when x"7AC" => DATA <= x"01";
            when x"7AD" => DATA <= x"7E";
            when x"7AE" => DATA <= x"F8";
            when x"7AF" => DATA <= x"F5";
            when x"7B0" => DATA <= x"7E";
            when x"7B1" => DATA <= x"F9";
            when x"7B2" => DATA <= x"4D";
            when x"7B3" => DATA <= x"7E";
            when x"7B4" => DATA <= x"F9";
            when x"7B5" => DATA <= x"1C";
            when x"7B6" => DATA <= x"7E";
            when x"7B7" => DATA <= x"F9";
            when x"7B8" => DATA <= x"4D";
            when x"7B9" => DATA <= x"7E";
            when x"7BA" => DATA <= x"F8";
            when x"7BB" => DATA <= x"67";
            when x"7BC" => DATA <= x"7E";
            when x"7BD" => DATA <= x"FD";
            when x"7BE" => DATA <= x"3F";
            when x"7BF" => DATA <= x"7E";
            when x"7C0" => DATA <= x"F8";
            when x"7C1" => DATA <= x"C3";
            when x"7C2" => DATA <= x"7E";
            when x"7C3" => DATA <= x"F9";
            when x"7C4" => DATA <= x"4D";
            when x"7C5" => DATA <= x"7E";
            when x"7C6" => DATA <= x"F9";
            when x"7C7" => DATA <= x"24";
            when x"7C8" => DATA <= x"7E";
            when x"7C9" => DATA <= x"F9";
            when x"7CA" => DATA <= x"4D";
            when x"7CB" => DATA <= x"7E";
            when x"7CC" => DATA <= x"F9";
            when x"7CD" => DATA <= x"4D";
            when x"7CE" => DATA <= x"7E";
            when x"7CF" => DATA <= x"FB";
            when x"7D0" => DATA <= x"1D";
            when x"7D1" => DATA <= x"7E";
            when x"7D2" => DATA <= x"FB";
            when x"7D3" => DATA <= x"6E";
            when x"7D4" => DATA <= x"7E";
            when x"7D5" => DATA <= x"FA";
            when x"7D6" => DATA <= x"F4";
            when x"7D7" => DATA <= x"7E";
            when x"7D8" => DATA <= x"FB";
            when x"7D9" => DATA <= x"05";
            when x"7DA" => DATA <= x"7E";
            when x"7DB" => DATA <= x"FA";
            when x"7DC" => DATA <= x"CE";
            when x"7DD" => DATA <= x"7E";
            when x"7DE" => DATA <= x"FB";
            when x"7DF" => DATA <= x"40";
            when x"7E0" => DATA <= x"7E";
            when x"7E1" => DATA <= x"F9";
            when x"7E2" => DATA <= x"2D";
            when x"7E3" => DATA <= x"81";
            when x"7E4" => DATA <= x"0D";
            when x"7E5" => DATA <= x"26";
            when x"7E6" => DATA <= x"07";
            when x"7E7" => DATA <= x"86";
            when x"7E8" => DATA <= x"0A";
            when x"7E9" => DATA <= x"BD";
            when x"7EA" => DATA <= x"FF";
            when x"7EB" => DATA <= x"EE";
            when x"7EC" => DATA <= x"86";
            when x"7ED" => DATA <= x"0D";
            when x"7EE" => DATA <= x"7E";
            when x"7EF" => DATA <= x"FB";
            when x"7F0" => DATA <= x"B9";
            when x"7F1" => DATA <= x"7E";
            when x"7F2" => DATA <= x"FA";
            when x"7F3" => DATA <= x"11";
            when x"7F4" => DATA <= x"7E";
            when x"7F5" => DATA <= x"F9";
            when x"7F6" => DATA <= x"9E";
            when x"7F7" => DATA <= x"7E";
            when x"7F8" => DATA <= x"F9";
            when x"7F9" => DATA <= x"3E";
            when x"7FA" => DATA <= x"F8";
            when x"7FB" => DATA <= x"A7";
            when x"7FC" => DATA <= x"F9";
            when x"7FD" => DATA <= x"4D";
            when x"7FE" => DATA <= x"F8";
            when x"7FF" => DATA <= x"2D";
            when others => DATA <= (others => '0');
        end case;
    end process;
end RTL;
